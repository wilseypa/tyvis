use std.textio.all;

entity ISCAS85_5 is 
	 generic (tpd_hl : time := 1 fs;
	          tpd_lh : time := 1 fs);
end;

architecture DEMO of ISCAS85_5 is

  signal  INP : bit_vector(0 to 32);
  signal  OUTP : bit_vector(0 to 24);
  signal  H : bit ;

 signal INTERP0 : bit := '0';
 signal INTERP1 : bit := '0';
 signal INTERP2 : bit := '0';
 signal INTERP3 : bit := '0';
 signal INTERP4 : bit := '0';
 signal INTERP5 : bit := '0';
 signal INTERP6 : bit := '0';
 signal INTERP7 : bit := '0';
 signal INTERP8 : bit := '0';
 signal INTERP9 : bit := '0';
 signal INTERP10 : bit := '0';
 signal INTERP11 : bit := '0';
 signal INTERP12 : bit := '0';
 signal INTERP13 : bit := '0';
 signal INTERP14 : bit := '0';
 signal INTERP15 : bit := '0';
 signal INTERP16 : bit := '0';
 signal INTERP17 : bit := '0';
 signal INTERP18 : bit := '0';
 signal INTERP19 : bit := '0';
 signal INTERP20 : bit := '0';
 signal INTERP21 : bit := '0';
 signal INTERP22 : bit := '0';
 signal INTERP23 : bit := '0';
 signal INTERP24 : bit := '0';
 signal INTERP25 : bit := '0';
 signal INTERP26 : bit := '0';
 signal INTERP27 : bit := '0';
 signal INTERP28 : bit := '0';
 signal INTERP29 : bit := '0';
 signal INTERP30 : bit := '0';
 signal INTERP31 : bit := '0';
 signal INTERP32 : bit := '0';
 signal INTERP33 : bit := '0';
 signal INTERP34 : bit := '0';
 signal INTERP35 : bit := '0';
 signal INTERP36 : bit := '0';
 signal INTERP37 : bit := '0';
 signal INTERP38 : bit := '0';
 signal INTERP39 : bit := '0';
 signal INTERP40 : bit := '0';
 signal INTERP41 : bit := '0';
 signal INTERP42 : bit := '0';
 signal INTERP43 : bit := '0';
 signal INTERP44 : bit := '0';
 signal INTERP45 : bit := '0';
 signal INTERP46 : bit := '0';
 signal INTERP47 : bit := '0';
 signal INTERP48 : bit := '0';
 signal INTERP49 : bit := '0';
 signal INTERP50 : bit := '0';
 signal INTERP51 : bit := '0';
 signal INTERP52 : bit := '0';
 signal INTERP53 : bit := '0';
 signal INTERP54 : bit := '0';
 signal INTERP55 : bit := '0';
 signal INTERP56 : bit := '0';
 signal INTERP57 : bit := '0';
 signal INTERP58 : bit := '0';
 signal INTERP59 : bit := '0';
 signal INTERP60 : bit := '0';
 signal INTERP61 : bit := '0';
 signal INTERP62 : bit := '0';
 signal INTERP63 : bit := '0';
 signal INTERP64 : bit := '0';
 signal INTERP65 : bit := '0';
 signal INTERP66 : bit := '0';
 signal INTERP67 : bit := '0';
 signal INTERP68 : bit := '0';
 signal INTERP69 : bit := '0';
 signal INTERP70 : bit := '0';
 signal INTERP71 : bit := '0';
 signal INTERP72 : bit := '0';
 signal INTERP73 : bit := '0';
 signal INTERP74 : bit := '0';
 signal INTERP75 : bit := '0';
 signal INTERP76 : bit := '0';
 signal INTERP77 : bit := '0';
 signal INTERP78 : bit := '0';
 signal INTERP79 : bit := '0';
 signal INTERP80 : bit := '0';
 signal INTERP81 : bit := '0';
 signal INTERP82 : bit := '0';
 signal INTERP83 : bit := '0';
 signal INTERP84 : bit := '0';
 signal INTERP85 : bit := '0';
 signal INTERP86 : bit := '0';
 signal INTERP87 : bit := '0';
 signal INTERP88 : bit := '0';
 signal INTERP89 : bit := '0';
 signal INTERP90 : bit := '0';
 signal INTERP91 : bit := '0';
 signal INTERP92 : bit := '0';
 signal INTERP93 : bit := '0';
 signal INTERP94 : bit := '0';
 signal INTERP95 : bit := '0';
 signal INTERP96 : bit := '0';
 signal INTERP97 : bit := '0';
 signal INTERP98 : bit := '0';
 signal INTERP99 : bit := '0';
 signal INTERP100 : bit := '0';
 signal INTERP101 : bit := '0';
 signal INTERP102 : bit := '0';
 signal INTERP103 : bit := '0';
 signal INTERP104 : bit := '0';
 signal INTERP105 : bit := '0';
 signal INTERP106 : bit := '0';
 signal INTERP107 : bit := '0';
 signal INTERP108 : bit := '0';
 signal INTERP109 : bit := '0';
 signal INTERP110 : bit := '0';
 signal INTERP111 : bit := '0';
 signal INTERP112 : bit := '0';
 signal INTERP113 : bit := '0';
 signal INTERP114 : bit := '0';
 signal INTERP115 : bit := '0';
 signal INTERP116 : bit := '0';
 signal INTERP117 : bit := '0';
 signal INTERP118 : bit := '0';
 signal INTERP119 : bit := '0';
 signal INTERP120 : bit := '0';
 signal INTERP121 : bit := '0';
 signal INTERP122 : bit := '0';
 signal INTERP123 : bit := '0';
 signal INTERP124 : bit := '0';
 signal INTERP125 : bit := '0';
 signal INTERP126 : bit := '0';
 signal INTERP127 : bit := '0';
 signal INTERP128 : bit := '0';
 signal INTERP129 : bit := '0';
 signal INTERP130 : bit := '0';
 signal INTERP131 : bit := '0';
 signal INTERP132 : bit := '0';
 signal INTERP133 : bit := '0';
 signal INTERP134 : bit := '0';
 signal INTERP135 : bit := '0';
 signal INTERP136 : bit := '0';
 signal INTERP137 : bit := '0';
 signal INTERP138 : bit := '0';
 signal INTERP139 : bit := '0';
 signal INTERP140 : bit := '0';
 signal INTERP141 : bit := '0';
 signal INTERP142 : bit := '0';
 signal INTERP143 : bit := '0';
 signal INTERP144 : bit := '0';
 signal INTERP145 : bit := '0';
 signal INTERP146 : bit := '0';
 signal INTERP147 : bit := '0';
 signal INTERP148 : bit := '0';
 signal INTERP149 : bit := '0';
 signal INTERP150 : bit := '0';
 signal INTERP151 : bit := '0';
 signal INTERP152 : bit := '0';
 signal INTERP153 : bit := '0';
 signal INTERP154 : bit := '0';
 signal INTERP155 : bit := '0';
 signal INTERP156 : bit := '0';
 signal INTERP157 : bit := '0';
 signal INTERP158 : bit := '0';
 signal INTERP159 : bit := '0';
 signal INTERP160 : bit := '0';
 signal INTERP161 : bit := '0';
 signal INTERP162 : bit := '0';
 signal INTERP163 : bit := '0';
 signal INTERP164 : bit := '0';
 signal INTERP165 : bit := '0';
 signal INTERP166 : bit := '0';
 signal INTERP167 : bit := '0';
 signal INTERP168 : bit := '0';
 signal INTERP169 : bit := '0';
 signal INTERP170 : bit := '0';
 signal INTERP171 : bit := '0';
 signal INTERP172 : bit := '0';
 signal INTERP173 : bit := '0';
 signal INTERP174 : bit := '0';
 signal INTERP175 : bit := '0';
 signal INTERP176 : bit := '0';
 signal INTERP177 : bit := '0';
 signal INTERP178 : bit := '0';
 signal INTERP179 : bit := '0';
 signal INTERP180 : bit := '0';
 signal INTERP181 : bit := '0';
 signal INTERP182 : bit := '0';
 signal INTERP183 : bit := '0';
 signal INTERP184 : bit := '0';
 signal INTERP185 : bit := '0';
 signal INTERP186 : bit := '0';
 signal INTERP187 : bit := '0';
 signal INTERP188 : bit := '0';
 signal INTERP189 : bit := '0';
 signal INTERP190 : bit := '0';
 signal INTERP191 : bit := '0';
 signal INTERP192 : bit := '0';
 signal INTERP193 : bit := '0';
 signal INTERP194 : bit := '0';
 signal INTERP195 : bit := '0';
 signal INTERP196 : bit := '0';
 signal INTERP197 : bit := '0';
 signal INTERP198 : bit := '0';
 signal INTERP199 : bit := '0';
 signal INTERP200 : bit := '0';
 signal INTERP201 : bit := '0';
 signal INTERP202 : bit := '0';
 signal INTERP203 : bit := '0';
 signal INTERP204 : bit := '0';
 signal INTERP205 : bit := '0';
 signal INTERP206 : bit := '0';
 signal INTERP207 : bit := '0';
 signal INTERP208 : bit := '0';
 signal INTERP209 : bit := '0';
 signal INTERP210 : bit := '0';
 signal INTERP211 : bit := '0';
 signal INTERP212 : bit := '0';
 signal INTERP213 : bit := '0';
 signal INTERP214 : bit := '0';
 signal INTERP215 : bit := '0';
 signal INTERP216 : bit := '0';
 signal INTERP217 : bit := '0';
 signal INTERP218 : bit := '0';
 signal INTERP219 : bit := '0';
 signal INTERP220 : bit := '0';
 signal INTERP221 : bit := '0';
 signal INTERP222 : bit := '0';
 signal INTERP223 : bit := '0';
 signal INTERP224 : bit := '0';
 signal INTERP225 : bit := '0';
 signal INTERP226 : bit := '0';
 signal INTERP227 : bit := '0';
 signal INTERP228 : bit := '0';
 signal INTERP229 : bit := '0';
 signal INTERP230 : bit := '0';
 signal INTERP231 : bit := '0';
 signal INTERP232 : bit := '0';
 signal INTERP233 : bit := '0';
 signal INTERP234 : bit := '0';
 signal INTERP235 : bit := '0';
 signal INTERP236 : bit := '0';
 signal INTERP237 : bit := '0';
 signal INTERP238 : bit := '0';
 signal INTERP239 : bit := '0';
 signal INTERP240 : bit := '0';
 signal INTERP241 : bit := '0';
 signal INTERP242 : bit := '0';
 signal INTERP243 : bit := '0';
 signal INTERP244 : bit := '0';
 signal INTERP245 : bit := '0';
 signal INTERP246 : bit := '0';
 signal INTERP247 : bit := '0';
 signal INTERP248 : bit := '0';
 signal INTERP249 : bit := '0';
 signal INTERP250 : bit := '0';
 signal INTERP251 : bit := '0';
 signal INTERP252 : bit := '0';
 signal INTERP253 : bit := '0';
 signal INTERP254 : bit := '0';
 signal INTERP255 : bit := '0';
 signal INTERP256 : bit := '0';
 signal INTERP257 : bit := '0';
 signal INTERP258 : bit := '0';
 signal INTERP259 : bit := '0';
 signal INTERP260 : bit := '0';
 signal INTERP261 : bit := '0';
 signal INTERP262 : bit := '0';
 signal INTERP263 : bit := '0';
 signal INTERP264 : bit := '0';
 signal INTERP265 : bit := '0';
 signal INTERP266 : bit := '0';
 signal INTERP267 : bit := '0';
 signal INTERP268 : bit := '0';
 signal INTERP269 : bit := '0';
 signal INTERP270 : bit := '0';
 signal INTERP271 : bit := '0';
 signal INTERP272 : bit := '0';
 signal INTERP273 : bit := '0';
 signal INTERP274 : bit := '0';
 signal INTERP275 : bit := '0';
 signal INTERP276 : bit := '0';
 signal INTERP277 : bit := '0';
 signal INTERP278 : bit := '0';
 signal INTERP279 : bit := '0';
 signal INTERP280 : bit := '0';
 signal INTERP281 : bit := '0';
 signal INTERP282 : bit := '0';
 signal INTERP283 : bit := '0';
 signal INTERP284 : bit := '0';
 signal INTERP285 : bit := '0';
 signal INTERP286 : bit := '0';
 signal INTERP287 : bit := '0';
 signal INTERP288 : bit := '0';
 signal INTERP289 : bit := '0';
 signal INTERP290 : bit := '0';
 signal INTERP291 : bit := '0';
 signal INTERP292 : bit := '0';
 signal INTERP293 : bit := '0';
 signal INTERP294 : bit := '0';
 signal INTERP295 : bit := '0';
 signal INTERP296 : bit := '0';
 signal INTERP297 : bit := '0';
 signal INTERP298 : bit := '0';
 signal INTERP299 : bit := '0';
 signal INTERP300 : bit := '0';
 signal INTERP301 : bit := '0';
 signal INTERP302 : bit := '0';
 signal INTERP303 : bit := '0';
 signal INTERP304 : bit := '0';
 signal INTERP305 : bit := '0';
 signal INTERP306 : bit := '0';
 signal INTERP307 : bit := '0';
 signal INTERP308 : bit := '0';
 signal INTERP309 : bit := '0';
 signal INTERP310 : bit := '0';
 signal INTERP311 : bit := '0';
 signal INTERP312 : bit := '0';
 signal INTERP313 : bit := '0';
 signal INTERP314 : bit := '0';
 signal INTERP315 : bit := '0';
 signal INTERP316 : bit := '0';
 signal INTERP317 : bit := '0';
 signal INTERP318 : bit := '0';
 signal INTERP319 : bit := '0';
 signal INTERP320 : bit := '0';
 signal INTERP321 : bit := '0';
 signal INTERP322 : bit := '0';
 signal INTERP323 : bit := '0';
 signal INTERP324 : bit := '0';
 signal INTERP325 : bit := '0';
 signal INTERP326 : bit := '0';
 signal INTERP327 : bit := '0';
 signal INTERP328 : bit := '0';
 signal INTERP329 : bit := '0';
 signal INTERP330 : bit := '0';
 signal INTERP331 : bit := '0';
 signal INTERP332 : bit := '0';
 signal INTERP333 : bit := '0';
 signal INTERP334 : bit := '0';
 signal INTERP335 : bit := '0';
 signal INTERP336 : bit := '0';
 signal INTERP337 : bit := '0';
 signal INTERP338 : bit := '0';
 signal INTERP339 : bit := '0';
 signal INTERP340 : bit := '0';
 signal INTERP341 : bit := '0';
 signal INTERP342 : bit := '0';
 signal INTERP343 : bit := '0';
 signal INTERP344 : bit := '0';
 signal INTERP345 : bit := '0';
 signal INTERP346 : bit := '0';
 signal INTERP347 : bit := '0';
 signal INTERP348 : bit := '0';
 signal INTERP349 : bit := '0';
 signal INTERP350 : bit := '0';
 signal INTERP351 : bit := '0';
 signal INTERP352 : bit := '0';
 signal INTERP353 : bit := '0';
 signal INTERP354 : bit := '0';
 signal INTERP355 : bit := '0';
 signal INTERP356 : bit := '0';
 signal INTERP357 : bit := '0';
 signal INTERP358 : bit := '0';
 signal INTERP359 : bit := '0';
 signal INTERP360 : bit := '0';
 signal INTERP361 : bit := '0';
 signal INTERP362 : bit := '0';
 signal INTERP363 : bit := '0';
 signal INTERP364 : bit := '0';
 signal INTERP365 : bit := '0';
 signal INTERP366 : bit := '0';
 signal INTERP367 : bit := '0';
 signal INTERP368 : bit := '0';
 signal INTERP369 : bit := '0';
 signal INTERP370 : bit := '0';
 signal INTERP371 : bit := '0';
 signal INTERP372 : bit := '0';
 signal INTERP373 : bit := '0';
 signal INTERP374 : bit := '0';
 signal INTERP375 : bit := '0';
 signal INTERP376 : bit := '0';
 signal INTERP377 : bit := '0';
 signal INTERP378 : bit := '0';
 signal INTERP379 : bit := '0';
 signal INTERP380 : bit := '0';
 signal INTERP381 : bit := '0';
 signal INTERP382 : bit := '0';
 signal INTERP383 : bit := '0';
 signal INTERP384 : bit := '0';
 signal INTERP385 : bit := '0';
 signal INTERP386 : bit := '0';
 signal INTERP387 : bit := '0';
 signal INTERP388 : bit := '0';
 signal INTERP389 : bit := '0';
 signal INTERP390 : bit := '0';
 signal INTERP391 : bit := '0';
 signal INTERP392 : bit := '0';
 signal INTERP393 : bit := '0';
 signal INTERP394 : bit := '0';
 signal INTERP395 : bit := '0';
 signal INTERP396 : bit := '0';
 signal INTERP397 : bit := '0';
 signal INTERP398 : bit := '0';
 signal INTERP399 : bit := '0';
 signal INTERP400 : bit := '0';
 signal INTERP401 : bit := '0';
 signal INTERP402 : bit := '0';
 signal INTERP403 : bit := '0';
 signal INTERP404 : bit := '0';
 signal INTERP405 : bit := '0';
 signal INTERP406 : bit := '0';
 signal INTERP407 : bit := '0';
 signal INTERP408 : bit := '0';
 signal INTERP409 : bit := '0';
 signal INTERP410 : bit := '0';
 signal INTERP411 : bit := '0';
 signal INTERP412 : bit := '0';
 signal INTERP413 : bit := '0';
 signal INTERP414 : bit := '0';
 signal INTERP415 : bit := '0';
 signal INTERP416 : bit := '0';
 signal INTERP417 : bit := '0';
 signal INTERP418 : bit := '0';
 signal INTERP419 : bit := '0';
 signal INTERP420 : bit := '0';
 signal INTERP421 : bit := '0';
 signal INTERP422 : bit := '0';
 signal INTERP423 : bit := '0';
 signal INTERP424 : bit := '0';
 signal INTERP425 : bit := '0';
 signal INTERP426 : bit := '0';
 signal INTERP427 : bit := '0';
 signal INTERP428 : bit := '0';
 signal INTERP429 : bit := '0';
 signal INTERP430 : bit := '0';
 signal INTERP431 : bit := '0';
 signal INTERP432 : bit := '0';
 signal INTERP433 : bit := '0';
 signal INTERP434 : bit := '0';
 signal INTERP435 : bit := '0';
 signal INTERP436 : bit := '0';
 signal INTERP437 : bit := '0';
 signal INTERP438 : bit := '0';
 signal INTERP439 : bit := '0';
 signal INTERP440 : bit := '0';
 signal INTERP441 : bit := '0';
 signal INTERP442 : bit := '0';
 signal INTERP443 : bit := '0';
 signal INTERP444 : bit := '0';
 signal INTERP445 : bit := '0';
 signal INTERP446 : bit := '0';
 signal INTERP447 : bit := '0';
 signal INTERP448 : bit := '0';
 signal INTERP449 : bit := '0';
 signal INTERP450 : bit := '0';
 signal INTERP451 : bit := '0';
 signal INTERP452 : bit := '0';
 signal INTERP453 : bit := '0';
 signal INTERP454 : bit := '0';
 signal INTERP455 : bit := '0';
 signal INTERP456 : bit := '0';
 signal INTERP457 : bit := '0';
 signal INTERP458 : bit := '0';
 signal INTERP459 : bit := '0';
 signal INTERP460 : bit := '0';
 signal INTERP461 : bit := '0';
 signal INTERP462 : bit := '0';
 signal INTERP463 : bit := '0';
 signal INTERP464 : bit := '0';
 signal INTERP465 : bit := '0';
 signal INTERP466 : bit := '0';
 signal INTERP467 : bit := '0';
 signal INTERP468 : bit := '0';
 signal INTERP469 : bit := '0';
 signal INTERP470 : bit := '0';
 signal INTERP471 : bit := '0';
 signal INTERP472 : bit := '0';
 signal INTERP473 : bit := '0';
 signal INTERP474 : bit := '0';
 signal INTERP475 : bit := '0';
 signal INTERP476 : bit := '0';
 signal INTERP477 : bit := '0';
 signal INTERP478 : bit := '0';
 signal INTERP479 : bit := '0';
 signal INTERP480 : bit := '0';
 signal INTERP481 : bit := '0';
 signal INTERP482 : bit := '0';
 signal INTERP483 : bit := '0';
 signal INTERP484 : bit := '0';
 signal INTERP485 : bit := '0';
 signal INTERP486 : bit := '0';
 signal INTERP487 : bit := '0';
 signal INTERP488 : bit := '0';
 signal INTERP489 : bit := '0';
 signal INTERP490 : bit := '0';
 signal INTERP491 : bit := '0';
 signal INTERP492 : bit := '0';
 signal INTERP493 : bit := '0';
 signal INTERP494 : bit := '0';
 signal INTERP495 : bit := '0';
 signal INTERP496 : bit := '0';
 signal INTERP497 : bit := '0';
 signal INTERP498 : bit := '0';
 signal INTERP499 : bit := '0';
 signal INTERP500 : bit := '0';
 signal INTERP501 : bit := '0';
 signal INTERP502 : bit := '0';
 signal INTERP503 : bit := '0';
 signal INTERP504 : bit := '0';
 signal INTERP505 : bit := '0';
 signal INTERP506 : bit := '0';
 signal INTERP507 : bit := '0';
 signal INTERP508 : bit := '0';
 signal INTERP509 : bit := '0';
 signal INTERP510 : bit := '0';
 signal INTERP511 : bit := '0';
 signal INTERP512 : bit := '0';
 signal INTERP513 : bit := '0';
 signal INTERP514 : bit := '0';
 signal INTERP515 : bit := '0';
 signal INTERP516 : bit := '0';
 signal INTERP517 : bit := '0';
 signal INTERP518 : bit := '0';
 signal INTERP519 : bit := '0';
 signal INTERP520 : bit := '0';
 signal INTERP521 : bit := '0';
 signal INTERP522 : bit := '0';
 signal INTERP523 : bit := '0';
 signal INTERP524 : bit := '0';
 signal INTERP525 : bit := '0';
 signal INTERP526 : bit := '0';
 signal INTERP527 : bit := '0';
 signal INTERP528 : bit := '0';
 signal INTERP529 : bit := '0';
 signal INTERP530 : bit := '0';
 signal INTERP531 : bit := '0';
 signal INTERP532 : bit := '0';
 signal INTERP533 : bit := '0';
 signal INTERP534 : bit := '0';
 signal INTERP535 : bit := '0';
 signal INTERP536 : bit := '0';
 signal INTERP537 : bit := '0';
 signal INTERP538 : bit := '0';
 signal INTERP539 : bit := '0';
 signal INTERP540 : bit := '0';
 signal INTERP541 : bit := '0';
 signal INTERP542 : bit := '0';
 signal INTERP543 : bit := '0';
 signal INTERP544 : bit := '0';
 signal INTERP545 : bit := '0';
 signal INTERP546 : bit := '0';
 signal INTERP547 : bit := '0';
 signal INTERP548 : bit := '0';
 signal INTERP549 : bit := '0';
 signal INTERP550 : bit := '0';
 signal INTERP551 : bit := '0';
 signal INTERP552 : bit := '0';
 signal INTERP553 : bit := '0';
 signal INTERP554 : bit := '0';
 signal INTERP555 : bit := '0';
 signal INTERP556 : bit := '0';
 signal INTERP557 : bit := '0';
 signal INTERP558 : bit := '0';
 signal INTERP559 : bit := '0';
 signal INTERP560 : bit := '0';
 signal INTERP561 : bit := '0';
 signal INTERP562 : bit := '0';
 signal INTERP563 : bit := '0';
 signal INTERP564 : bit := '0';
 signal INTERP565 : bit := '0';
 signal INTERP566 : bit := '0';
 signal INTERP567 : bit := '0';
 signal INTERP568 : bit := '0';
 signal INTERP569 : bit := '0';
 signal INTERP570 : bit := '0';
 signal INTERP571 : bit := '0';
 signal INTERP572 : bit := '0';
 signal INTERP573 : bit := '0';
 signal INTERP574 : bit := '0';
 signal INTERP575 : bit := '0';
 signal INTERP576 : bit := '0';
 signal INTERP577 : bit := '0';
 signal INTERP578 : bit := '0';
 signal INTERP579 : bit := '0';
 signal INTERP580 : bit := '0';
 signal INTERP581 : bit := '0';
 signal INTERP582 : bit := '0';
 signal INTERP583 : bit := '0';
 signal INTERP584 : bit := '0';
 signal INTERP585 : bit := '0';
 signal INTERP586 : bit := '0';
 signal INTERP587 : bit := '0';
 signal INTERP588 : bit := '0';
 signal INTERP589 : bit := '0';
 signal INTERP590 : bit := '0';
 signal INTERP591 : bit := '0';
 signal INTERP592 : bit := '0';
 signal INTERP593 : bit := '0';
 signal INTERP594 : bit := '0';
 signal INTERP595 : bit := '0';
 signal INTERP596 : bit := '0';
 signal INTERP597 : bit := '0';
 signal INTERP598 : bit := '0';
 signal INTERP599 : bit := '0';
 signal INTERP600 : bit := '0';
 signal INTERP601 : bit := '0';
 signal INTERP602 : bit := '0';
 signal INTERP603 : bit := '0';
 signal INTERP604 : bit := '0';
 signal INTERP605 : bit := '0';
 signal INTERP606 : bit := '0';
 signal INTERP607 : bit := '0';
 signal INTERP608 : bit := '0';
 signal INTERP609 : bit := '0';
 signal INTERP610 : bit := '0';
 signal INTERP611 : bit := '0';
 signal INTERP612 : bit := '0';
 signal INTERP613 : bit := '0';
 signal INTERP614 : bit := '0';
 signal INTERP615 : bit := '0';
 signal INTERP616 : bit := '0';
 signal INTERP617 : bit := '0';
 signal INTERP618 : bit := '0';
 signal INTERP619 : bit := '0';
 signal INTERP620 : bit := '0';
 signal INTERP621 : bit := '0';
 signal INTERP622 : bit := '0';
 signal INTERP623 : bit := '0';
 signal INTERP624 : bit := '0';
 signal INTERP625 : bit := '0';
 signal INTERP626 : bit := '0';
 signal INTERP627 : bit := '0';
 signal INTERP628 : bit := '0';
 signal INTERP629 : bit := '0';
 signal INTERP630 : bit := '0';
 signal INTERP631 : bit := '0';
 signal INTERP632 : bit := '0';
 signal INTERP633 : bit := '0';
 signal INTERP634 : bit := '0';
 signal INTERP635 : bit := '0';
 signal INTERP636 : bit := '0';
 signal INTERP637 : bit := '0';
 signal INTERP638 : bit := '0';
 signal INTERP639 : bit := '0';
 signal INTERP640 : bit := '0';
 signal INTERP641 : bit := '0';
 signal INTERP642 : bit := '0';
 signal INTERP643 : bit := '0';
 signal INTERP644 : bit := '0';
 signal INTERP645 : bit := '0';
 signal INTERP646 : bit := '0';
 signal INTERP647 : bit := '0';
 signal INTERP648 : bit := '0';
 signal INTERP649 : bit := '0';
 signal INTERP650 : bit := '0';
 signal INTERP651 : bit := '0';
 signal INTERP652 : bit := '0';
 signal INTERP653 : bit := '0';
 signal INTERP654 : bit := '0';
 signal INTERP655 : bit := '0';
 signal INTERP656 : bit := '0';
 signal INTERP657 : bit := '0';
 signal INTERP658 : bit := '0';
 signal INTERP659 : bit := '0';
 signal INTERP660 : bit := '0';
 signal INTERP661 : bit := '0';
 signal INTERP662 : bit := '0';
 signal INTERP663 : bit := '0';
 signal INTERP664 : bit := '0';
 signal INTERP665 : bit := '0';
 signal INTERP666 : bit := '0';
 signal INTERP667 : bit := '0';
 signal INTERP668 : bit := '0';
 signal INTERP669 : bit := '0';
 signal INTERP670 : bit := '0';
 signal INTERP671 : bit := '0';
 signal INTERP672 : bit := '0';
 signal INTERP673 : bit := '0';
 signal INTERP674 : bit := '0';
 signal INTERP675 : bit := '0';
 signal INTERP676 : bit := '0';
 signal INTERP677 : bit := '0';
 signal INTERP678 : bit := '0';
 signal INTERP679 : bit := '0';
 signal INTERP680 : bit := '0';
 signal INTERP681 : bit := '0';
 signal INTERP682 : bit := '0';
 signal INTERP683 : bit := '0';
 signal INTERP684 : bit := '0';
 signal INTERP685 : bit := '0';
 signal INTERP686 : bit := '0';
 signal INTERP687 : bit := '0';
 signal INTERP688 : bit := '0';
 signal INTERP689 : bit := '0';
 signal INTERP690 : bit := '0';
 signal INTERP691 : bit := '0';
 signal INTERP692 : bit := '0';
 signal INTERP693 : bit := '0';
 signal INTERP694 : bit := '0';
 signal INTERP695 : bit := '0';
 signal INTERP696 : bit := '0';
 signal INTERP697 : bit := '0';
 signal INTERP698 : bit := '0';
 signal INTERP699 : bit := '0';
 signal INTERP700 : bit := '0';
 signal INTERP701 : bit := '0';
 signal INTERP702 : bit := '0';
 signal INTERP703 : bit := '0';
 signal INTERP704 : bit := '0';
 signal INTERP705 : bit := '0';
 signal INTERP706 : bit := '0';
 signal INTERP707 : bit := '0';
 signal INTERP708 : bit := '0';
 signal INTERP709 : bit := '0';
 signal INTERP710 : bit := '0';
 signal INTERP711 : bit := '0';
 signal INTERP712 : bit := '0';
 signal INTERP713 : bit := '0';
 signal INTERP714 : bit := '0';
 signal INTERP715 : bit := '0';
 signal INTERP716 : bit := '0';
 signal INTERP717 : bit := '0';
 signal INTERP718 : bit := '0';
 signal INTERP719 : bit := '0';
 signal INTERP720 : bit := '0';
 signal INTERP721 : bit := '0';
 signal INTERP722 : bit := '0';
 signal INTERP723 : bit := '0';
 signal INTERP724 : bit := '0';
 signal INTERP725 : bit := '0';
 signal INTERP726 : bit := '0';
 signal INTERP727 : bit := '0';
 signal INTERP728 : bit := '0';
 signal INTERP729 : bit := '0';
 signal INTERP730 : bit := '0';
 signal INTERP731 : bit := '0';
 signal INTERP732 : bit := '0';
 signal INTERP733 : bit := '0';
 signal INTERP734 : bit := '0';
 signal INTERP735 : bit := '0';
 signal INTERP736 : bit := '0';
 signal INTERP737 : bit := '0';
 signal INTERP738 : bit := '0';
 signal INTERP739 : bit := '0';
 signal INTERP740 : bit := '0';
 signal INTERP741 : bit := '0';
 signal INTERP742 : bit := '0';
 signal INTERP743 : bit := '0';
 signal INTERP744 : bit := '0';
 signal INTERP745 : bit := '0';
 signal INTERP746 : bit := '0';
 signal INTERP747 : bit := '0';
 signal INTERP748 : bit := '0';
 signal INTERP749 : bit := '0';
 signal INTERP750 : bit := '0';
 signal INTERP751 : bit := '0';
 signal INTERP752 : bit := '0';
 signal INTERP753 : bit := '0';
 signal INTERP754 : bit := '0';
 signal INTERP755 : bit := '0';
 signal INTERP756 : bit := '0';
 signal INTERP757 : bit := '0';
 signal INTERP758 : bit := '0';
 signal INTERP759 : bit := '0';
 signal INTERP760 : bit := '0';
 signal INTERP761 : bit := '0';
 signal INTERP762 : bit := '0';
 signal INTERP763 : bit := '0';
 signal INTERP764 : bit := '0';
 signal INTERP765 : bit := '0';
 signal INTERP766 : bit := '0';
 signal INTERP767 : bit := '0';
 signal INTERP768 : bit := '0';
 signal INTERP769 : bit := '0';
 signal INTERP770 : bit := '0';
 signal INTERP771 : bit := '0';
 signal INTERP772 : bit := '0';
 signal INTERP773 : bit := '0';
 signal INTERP774 : bit := '0';
 signal INTERP775 : bit := '0';
 signal INTERP776 : bit := '0';
 signal INTERP777 : bit := '0';
 signal INTERP778 : bit := '0';
 signal INTERP779 : bit := '0';
 signal INTERP780 : bit := '0';
 signal INTERP781 : bit := '0';
 signal INTERP782 : bit := '0';
 signal INTERP783 : bit := '0';
 signal INTERP784 : bit := '0';
 signal INTERP785 : bit := '0';
 signal INTERP786 : bit := '0';
 signal INTERP787 : bit := '0';
 signal INTERP788 : bit := '0';
 signal INTERP789 : bit := '0';
 signal INTERP790 : bit := '0';
 signal INTERP791 : bit := '0';
 signal INTERP792 : bit := '0';
 signal INTERP793 : bit := '0';
 signal INTERP794 : bit := '0';
 signal INTERP795 : bit := '0';
 signal INTERP796 : bit := '0';
 signal INTERP797 : bit := '0';
 signal INTERP798 : bit := '0';
 signal INTERP799 : bit := '0';
 signal INTERP800 : bit := '0';
 signal INTERP801 : bit := '0';
 signal INTERP802 : bit := '0';
 signal INTERP803 : bit := '0';
 signal INTERP804 : bit := '0';
 signal INTERP805 : bit := '0';
 signal INTERP806 : bit := '0';
 signal INTERP807 : bit := '0';
 signal INTERP808 : bit := '0';
 signal INTERP809 : bit := '0';
 signal INTERP810 : bit := '0';
 signal INTERP811 : bit := '0';
 signal INTERP812 : bit := '0';
 signal INTERP813 : bit := '0';
 signal INTERP814 : bit := '0';
 signal INTERP815 : bit := '0';
 signal INTERP816 : bit := '0';
 signal INTERP817 : bit := '0';
 signal INTERP818 : bit := '0';
 signal INTERP819 : bit := '0';
 signal INTERP820 : bit := '0';
 signal INTERP821 : bit := '0';
 signal INTERP822 : bit := '0';
 signal INTERP823 : bit := '0';
 signal INTERP824 : bit := '0';
 signal INTERP825 : bit := '0';
 signal INTERP826 : bit := '0';
 signal INTERP827 : bit := '0';
 signal INTERP828 : bit := '0';
 signal INTERP829 : bit := '0';
 signal INTERP830 : bit := '0';
 signal INTERP831 : bit := '0';
 signal INTERP832 : bit := '0';
 signal INTERP833 : bit := '0';
 signal INTERP834 : bit := '0';
 signal INTERP835 : bit := '0';
 signal INTERP836 : bit := '0';
 signal INTERP837 : bit := '0';
 signal INTERP838 : bit := '0';
 signal INTERP839 : bit := '0';
 signal INTERP840 : bit := '0';
 signal INTERP841 : bit := '0';
 signal INTERP842 : bit := '0';
 signal INTERP843 : bit := '0';
 signal INTERP844 : bit := '0';
 signal INTERP845 : bit := '0';
 signal INTERP846 : bit := '0';
 signal INTERP847 : bit := '0';
 signal INTERP848 : bit := '0';
 signal INTERP849 : bit := '0';
 signal INTERP850 : bit := '0';
 signal INTERP851 : bit := '0';
 signal INTERP852 : bit := '0';
 signal INTERP853 : bit := '0';
 signal INTERP854 : bit := '0';
 signal INTERP855 : bit := '0';
 signal INTERP856 : bit := '0';
 signal INTERP857 : bit := '0';
 signal INTERP858 : bit := '0';
 signal INTERP859 : bit := '0';
 signal INTERP860 : bit := '0';
 signal INTERP861 : bit := '0';
 signal INTERP862 : bit := '0';
 signal INTERP863 : bit := '0';
 signal INTERP864 : bit := '0';
 signal INTERP865 : bit := '0';
 signal INTERP866 : bit := '0';
 signal INTERP867 : bit := '0';
 signal INTERP868 : bit := '0';
 signal INTERP869 : bit := '0';
 signal INTERP870 : bit := '0';
 signal INTERP871 : bit := '0';
 signal INTERP872 : bit := '0';
 signal INTERP873 : bit := '0';
 signal INTERP874 : bit := '0';
 signal INTERP875 : bit := '0';
 signal INTERP876 : bit := '0';
 signal INTERP877 : bit := '0';
 signal INTERP878 : bit := '0';
 signal INTERP879 : bit := '0';
 signal INTERP880 : bit := '0';
 signal INTERP881 : bit := '0';
 signal INTERP882 : bit := '0';
 signal INTERP883 : bit := '0';
 signal INTERP884 : bit := '0';
 signal INTERP885 : bit := '0';
 signal INTERP886 : bit := '0';
 signal INTERP887 : bit := '0';
 signal INTERP888 : bit := '0';
 signal INTERP889 : bit := '0';
 signal INTERP890 : bit := '0';
 signal INTERP891 : bit := '0';
 signal INTERP892 : bit := '0';
 signal INTERP893 : bit := '0';
 signal INTERP894 : bit := '0';
 signal INTERP895 : bit := '0';
 signal INTERP896 : bit := '0';
 signal INTERP897 : bit := '0';
 signal INTERP898 : bit := '0';
 signal INTERP899 : bit := '0';
 signal INTERP900 : bit := '0';
 signal INTERP901 : bit := '0';
 signal INTERP902 : bit := '0';
 signal INTERP903 : bit := '0';
 signal INTERP904 : bit := '0';
 signal INTERP905 : bit := '0';
 signal INTERP906 : bit := '0';
 signal INTERP907 : bit := '0';
 signal INTERP908 : bit := '0';
 signal INTERP909 : bit := '0';
 signal INTERP910 : bit := '0';
 signal INTERP911 : bit := '0';
 signal INTERP912 : bit := '0';
 signal INTERP913 : bit := '0';
 signal INTERP914 : bit := '0';
 signal INTERP915 : bit := '0';
 signal INTERP916 : bit := '0';
 signal INTERP917 : bit := '0';
 signal INTERP918 : bit := '0';
 signal INTERP919 : bit := '0';
 signal INTERP920 : bit := '0';
 signal INTERP921 : bit := '0';
 signal INTERP922 : bit := '0';
 signal INTERP923 : bit := '0';
 signal INTERP924 : bit := '0';
 signal INTERP925 : bit := '0';
 signal INTERP926 : bit := '0';
 signal INTERP927 : bit := '0';
 signal INTERP928 : bit := '0';
 signal INTERP929 : bit := '0';
 signal INTERP930 : bit := '0';
 signal INTERP931 : bit := '0';
 signal INTERP932 : bit := '0';
 signal INTERP933 : bit := '0';
 signal INTERP934 : bit := '0';
 signal INTERP935 : bit := '0';
 signal INTERP936 : bit := '0';
 signal INTERP937 : bit := '0';
 signal INTERP938 : bit := '0';
 signal INTERP939 : bit := '0';
 signal INTERP940 : bit := '0';
 signal INTERP941 : bit := '0';
 signal INTERP942 : bit := '0';
 signal INTERP943 : bit := '0';
 signal INTERP944 : bit := '0';
 signal INTERP945 : bit := '0';
 signal INTERP946 : bit := '0';
 signal INTERP947 : bit := '0';
 signal INTERP948 : bit := '0';
 signal INTERP949 : bit := '0';
 signal INTERP950 : bit := '0';
 signal INTERP951 : bit := '0';
 signal INTERP952 : bit := '0';
 signal INTERP953 : bit := '0';
 signal INTERP954 : bit := '0';
 signal INTERP955 : bit := '0';
 signal INTERP956 : bit := '0';
 signal INTERP957 : bit := '0';
 signal INTERP958 : bit := '0';
 signal INTERP959 : bit := '0';
 signal INTERP960 : bit := '0';
 signal INTERP961 : bit := '0';
 signal INTERP962 : bit := '0';
 signal INTERP963 : bit := '0';
 signal INTERP964 : bit := '0';
 signal INTERP965 : bit := '0';
 signal INTERP966 : bit := '0';
 signal INTERP967 : bit := '0';
 signal INTERP968 : bit := '0';
 signal INTERP969 : bit := '0';
 signal INTERP970 : bit := '0';
 signal INTERP971 : bit := '0';
 signal INTERP972 : bit := '0';
 signal INTERP973 : bit := '0';
 signal INTERP974 : bit := '0';
 signal INTERP975 : bit := '0';
 signal INTERP976 : bit := '0';
 signal INTERP977 : bit := '0';
 signal INTERP978 : bit := '0';
 signal INTERP979 : bit := '0';
 signal INTERP980 : bit := '0';
 signal INTERP981 : bit := '0';
 signal INTERP982 : bit := '0';
 signal INTERP983 : bit := '0';
 signal INTERP984 : bit := '0';
 signal INTERP985 : bit := '0';
 signal INTERP986 : bit := '0';
 signal INTERP987 : bit := '0';
 signal INTERP988 : bit := '0';
 signal INTERP989 : bit := '0';
 signal INTERP990 : bit := '0';
 signal INTERP991 : bit := '0';
 signal INTERP992 : bit := '0';
 signal INTERP993 : bit := '0';
 signal INTERP994 : bit := '0';
 signal INTERP995 : bit := '0';
 signal INTERP996 : bit := '0';
 signal INTERP997 : bit := '0';
 signal INTERP998 : bit := '0';
 signal INTERP999 : bit := '0';
 signal INTERP1000 : bit := '0';
 signal INTERP1001 : bit := '0';
 signal INTERP1002 : bit := '0';
 signal INTERP1003 : bit := '0';
 signal INTERP1004 : bit := '0';
 signal INTERP1005 : bit := '0';
 signal INTERP1006 : bit := '0';
 signal INTERP1007 : bit := '0';
 signal INTERP1008 : bit := '0';
 signal INTERP1009 : bit := '0';
 signal INTERP1010 : bit := '0';
 signal INTERP1011 : bit := '0';
 signal INTERP1012 : bit := '0';
 signal INTERP1013 : bit := '0';
 signal INTERP1014 : bit := '0';
 signal INTERP1015 : bit := '0';
 signal INTERP1016 : bit := '0';
 signal INTERP1017 : bit := '0';
 signal INTERP1018 : bit := '0';
 signal INTERP1019 : bit := '0';
 signal INTERP1020 : bit := '0';
 signal INTERP1021 : bit := '0';
 signal INTERP1022 : bit := '0';
 signal INTERP1023 : bit := '0';
 signal INTERP1024 : bit := '0';
 signal INTERP1025 : bit := '0';
 signal INTERP1026 : bit := '0';
 signal INTERP1027 : bit := '0';
 signal INTERP1028 : bit := '0';
 signal INTERP1029 : bit := '0';
 signal INTERP1030 : bit := '0';
 signal INTERP1031 : bit := '0';
 signal INTERP1032 : bit := '0';
 signal INTERP1033 : bit := '0';
 signal INTERP1034 : bit := '0';
 signal INTERP1035 : bit := '0';
 signal INTERP1036 : bit := '0';
 signal OUTPI : bit_vector(OUTP'range):=(others=>'0') ;

BEGIN


      INV0 : process(INP(0))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(0));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP0 <= val after tpd_hl;
            when '1' =>
                INTERP0 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV1 : process(INP(1))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(1));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1 <= val after tpd_hl;
            when '1' =>
                INTERP1 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV2 : process(INP(2))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(2));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP2 <= val after tpd_hl;
            when '1' =>
                INTERP2 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV3 : process(INP(3))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(3));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP3 <= val after tpd_hl;
            when '1' =>
                INTERP3 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV4 : process(INP(4))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(4));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP4 <= val after tpd_hl;
            when '1' =>
                INTERP4 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV5 : process(INP(5))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(5));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP5 <= val after tpd_hl;
            when '1' =>
                INTERP5 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV6 : process(INP(6))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(6));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP6 <= val after tpd_hl;
            when '1' =>
                INTERP6 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV7 : process(INP(7))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(7));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP7 <= val after tpd_hl;
            when '1' =>
                INTERP7 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV8 : process(INP(8))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(8));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP8 <= val after tpd_hl;
            when '1' =>
                INTERP8 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV9 : process(INP(9))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(9));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP9 <= val after tpd_hl;
            when '1' =>
                INTERP9 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV10 : process(INP(10))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(10));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP10 <= val after tpd_hl;
            when '1' =>
                INTERP10 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV11 : process(INP(11))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(11));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP11 <= val after tpd_hl;
            when '1' =>
                INTERP11 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV12 : process(INP(12))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(12));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP12 <= val after tpd_hl;
            when '1' =>
                INTERP12 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV13 : process(INP(13))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(13));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP13 <= val after tpd_hl;
            when '1' =>
                INTERP13 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV14 : process(INP(14))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(14));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP14 <= val after tpd_hl;
            when '1' =>
                INTERP14 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV15 : process(INP(15))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(15));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP15 <= val after tpd_hl;
            when '1' =>
                INTERP15 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND0 : process(INP(20), INP(28))
        variable val,ex_value : bit := '0';
    begin
        val := not(INP(20) and INP(28));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP16 <= val after tpd_hl;
            when '1' =>
                INTERP16 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND1 : process(INP(21), INP(29))
        variable val,ex_value : bit := '0';
    begin
        val := not(INP(21) and INP(29));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP17 <= val after tpd_hl;
            when '1' =>
                INTERP17 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV16 : process(INP(23))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(23));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP18 <= val after tpd_hl;
            when '1' =>
                INTERP18 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV17 : process(INP(23))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(23));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP19 <= val after tpd_hl;
            when '1' =>
                INTERP19 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV18 : process(INP(24))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(24));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP20 <= val after tpd_hl;
            when '1' =>
                INTERP20 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV19 : process(INP(25))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(25));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP21 <= val after tpd_hl;
            when '1' =>
                INTERP21 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV20 : process(INP(26))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(26));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP22 <= val after tpd_hl;
            when '1' =>
                INTERP22 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV21 : process(INP(27))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(27));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP23 <= val after tpd_hl;
            when '1' =>
                INTERP23 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV22 : process(INP(32))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(32));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP24 <= val after tpd_hl;
            when '1' =>
                INTERP24 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV23 : process(INP(32))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(32));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP25 <= val after tpd_hl;
            when '1' =>
                INTERP25 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV24 : process(INP(28))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(28));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP26 <= val after tpd_hl;
            when '1' =>
                INTERP26 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV25 : process(INP(29))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(29));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP27 <= val after tpd_hl;
            when '1' =>
                INTERP27 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV26 : process(INP(30))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(30));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP28 <= val after tpd_hl;
            when '1' =>
                INTERP28 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV27 : process(INP(30))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(30));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP29 <= val after tpd_hl;
            when '1' =>
                INTERP29 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV28 : process(INP(31))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(31));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP30 <= val after tpd_hl;
            when '1' =>
                INTERP30 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV29 : process(INP(31))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(31));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP31 <= val after tpd_hl;
            when '1' =>
                INTERP31 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV30 : process(INP(32))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(32));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP32 <= val after tpd_hl;
            when '1' =>
                INTERP32 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV31 : process(INP(32))
        variable val,ex_value : bit := '0';

    begin
        val := not(INP(32));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP33 <= val after tpd_hl;
            when '1' =>
                INTERP33 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV32 : process(INTERP35)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP35);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP34 <= val after tpd_hl;
            when '1' =>
                INTERP34 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV33 : process(INTERP37)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP37);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP36 <= val after tpd_hl;
            when '1' =>
                INTERP36 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV34 : process(INTERP39)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP39);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP38 <= val after tpd_hl;
            when '1' =>
                INTERP38 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV35 : process(INTERP41)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP41);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP40 <= val after tpd_hl;
            when '1' =>
                INTERP40 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV36 : process(INTERP43)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP43);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP42 <= val after tpd_hl;
            when '1' =>
                INTERP42 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV37 : process(INTERP45)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP45);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP44 <= val after tpd_hl;
            when '1' =>
                INTERP44 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV38 : process(INTERP47)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP47);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP46 <= val after tpd_hl;
            when '1' =>
                INTERP46 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV39 : process(INTERP49)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP49);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP48 <= val after tpd_hl;
            when '1' =>
                INTERP48 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV40 : process(INTERP51)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP51);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP50 <= val after tpd_hl;
            when '1' =>
                INTERP50 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV41 : process(INTERP53)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP53);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP52 <= val after tpd_hl;
            when '1' =>
                INTERP52 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV42 : process(INTERP55)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP55);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP54 <= val after tpd_hl;
            when '1' =>
                INTERP54 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV43 : process(INTERP57)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP57);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP56 <= val after tpd_hl;
            when '1' =>
                INTERP56 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV44 : process(INTERP59)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP59);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP58 <= val after tpd_hl;
            when '1' =>
                INTERP58 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV45 : process(INTERP61)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP61);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP60 <= val after tpd_hl;
            when '1' =>
                INTERP60 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV46 : process(INTERP63)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP63);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP62 <= val after tpd_hl;
            when '1' =>
                INTERP62 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV47 : process(INTERP65)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP65);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP64 <= val after tpd_hl;
            when '1' =>
                INTERP64 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND2 : process(INTERP30, INTERP67)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP30 and INTERP67);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP66 <= val after tpd_hl;
            when '1' =>
                INTERP66 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND3 : process(INTERP30, INTERP69)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP30 and INTERP69);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP68 <= val after tpd_hl;
            when '1' =>
                INTERP68 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND4 : process(INTERP30, INTERP71)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP30 and INTERP71);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP70 <= val after tpd_hl;
            when '1' =>
                INTERP70 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND5 : process(INTERP30, INTERP73)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP30 and INTERP73);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP72 <= val after tpd_hl;
            when '1' =>
                INTERP72 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND6 : process(INTERP30, INTERP75)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP30 and INTERP75);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP74 <= val after tpd_hl;
            when '1' =>
                INTERP74 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND7 : process(INTERP30, INTERP77)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP30 and INTERP77);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP76 <= val after tpd_hl;
            when '1' =>
                INTERP76 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND0 : process(INP(20), INTERP32)
        variable val,ex_value : bit := '0';
    begin
        val := INP(20) and INTERP32;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP78 <= val after tpd_hl;
            when '1' =>
                INTERP78 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND1 : process(INP(21), INTERP32)
        variable val,ex_value : bit := '0';
    begin
        val := INP(21) and INTERP32;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP79 <= val after tpd_hl;
            when '1' =>
                INTERP79 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND8 : process(INTERP82, INTERP26)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP82 and INTERP26);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP81 <= val after tpd_hl;
            when '1' =>
                INTERP81 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND9 : process(INTERP84, INTERP27)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP84 and INTERP27);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP83 <= val after tpd_hl;
            when '1' =>
                INTERP83 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND10 : process(INTERP86, INP(23))
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP86 and INP(23));

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP85 <= val after tpd_hl;
            when '1' =>
                INTERP85 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND11 : process(INTERP88, INTERP29)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP88 and INTERP29);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP87 <= val after tpd_hl;
            when '1' =>
                INTERP87 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND12 : process(INTERP19, INTERP29)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP19 and INTERP29);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP89 <= val after tpd_hl;
            when '1' =>
                INTERP89 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND5 : process(INTERP16, INTERP95)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP16 and INTERP95;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP94 <= val after tpd_hl;
            when '1' =>
                INTERP94 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND6 : process(INTERP17, INTERP97)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP17 and INTERP97;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP96 <= val after tpd_hl;
            when '1' =>
                INTERP96 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV48 : process(INTERP94)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP94);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP99 <= val after tpd_hl;
            when '1' =>
                INTERP99 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV49 : process(INTERP96)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP96);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP100 <= val after tpd_hl;
            when '1' =>
                INTERP100 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV50 : process(INTERP102)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP102);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP101 <= val after tpd_hl;
            when '1' =>
                INTERP101 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV51 : process(INTERP104)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP104);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP103 <= val after tpd_hl;
            when '1' =>
                INTERP103 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV52 : process(INTERP106)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP106);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP105 <= val after tpd_hl;
            when '1' =>
                INTERP105 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV53 : process(INTERP108)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP108);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP107 <= val after tpd_hl;
            when '1' =>
                INTERP107 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV54 : process(INTERP110)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP110);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP109 <= val after tpd_hl;
            when '1' =>
                INTERP109 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV55 : process(INTERP90)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP90);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP111 <= val after tpd_hl;
            when '1' =>
                INTERP111 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV56 : process(INTERP113)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP113);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP112 <= val after tpd_hl;
            when '1' =>
                INTERP112 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV57 : process(INTERP115)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP115);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP114 <= val after tpd_hl;
            when '1' =>
                INTERP114 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV58 : process(INTERP92)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP92);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP116 <= val after tpd_hl;
            when '1' =>
                INTERP116 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND8 : process(INP(16), INTERP89)
        variable val,ex_value : bit := '0';
    begin
        val := INP(16) and INTERP89;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP117 <= val after tpd_hl;
            when '1' =>
                INTERP117 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND9 : process(INP(18), INTERP87)
        variable val,ex_value : bit := '0';
    begin
        val := INP(18) and INTERP87;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP118 <= val after tpd_hl;
            when '1' =>
                INTERP118 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND13 : process(INP(17), INTERP89)
        variable val,ex_value : bit := '0';
    begin
        val := not(INP(17) and INTERP89);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP119 <= val after tpd_hl;
            when '1' =>
                INTERP119 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND14 : process(INP(19), INTERP87)
        variable val,ex_value : bit := '0';
    begin
        val := not(INP(19) and INTERP87);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP120 <= val after tpd_hl;
            when '1' =>
                INTERP120 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND15 : process(INP(16), INTERP89)
        variable val,ex_value : bit := '0';
    begin
        val := not(INP(16) and INTERP89);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP121 <= val after tpd_hl;
            when '1' =>
                INTERP121 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND16 : process(INP(18), INTERP87)
        variable val,ex_value : bit := '0';
    begin
        val := not(INP(18) and INTERP87);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP122 <= val after tpd_hl;
            when '1' =>
                INTERP122 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV59 : process(INTERP124)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP124);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP123 <= val after tpd_hl;
            when '1' =>
                INTERP123 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV60 : process(INTERP126)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP126);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP125 <= val after tpd_hl;
            when '1' =>
                INTERP125 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV61 : process(INTERP128)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP128);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP127 <= val after tpd_hl;
            when '1' =>
                INTERP127 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV62 : process(INTERP130)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP130);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP129 <= val after tpd_hl;
            when '1' =>
                INTERP129 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV63 : process(INTERP132)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP132);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP131 <= val after tpd_hl;
            when '1' =>
                INTERP131 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV64 : process(INTERP134)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP134);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP133 <= val after tpd_hl;
            when '1' =>
                INTERP133 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV65 : process(INTERP136)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP136);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP135 <= val after tpd_hl;
            when '1' =>
                INTERP135 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV66 : process(INTERP138)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP138);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP137 <= val after tpd_hl;
            when '1' =>
                INTERP137 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;

  NAND17 :
 INTERP139 <= not(INTERP26 and INTERP140 and INTERP141 and INTERP85) after tpd_hl;

  NAND18 :
 INTERP142 <= not(INTERP27 and INTERP143 and INTERP144 and INTERP85) after tpd_hl;

  NAND19 :
 INTERP145 <= not(INTERP146 and INTERP33 and INTERP85) after tpd_hl;


      INV67 : process(INTERP150)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP150);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP149 <= val after tpd_hl;
            when '1' =>
                INTERP149 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV68 : process(INTERP152)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP152);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP151 <= val after tpd_hl;
            when '1' =>
                INTERP151 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV69 : process(INTERP154)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP154);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP153 <= val after tpd_hl;
            when '1' =>
                INTERP153 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV70 : process(INTERP156)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP156);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP155 <= val after tpd_hl;
            when '1' =>
                INTERP155 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV71 : process(INTERP158)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP158);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP157 <= val after tpd_hl;
            when '1' =>
                INTERP157 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV72 : process(INTERP160)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP160);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP159 <= val after tpd_hl;
            when '1' =>
                INTERP159 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV73 : process(INTERP162)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP162);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP161 <= val after tpd_hl;
            when '1' =>
                INTERP161 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV74 : process(INTERP164)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP164);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP163 <= val after tpd_hl;
            when '1' =>
                INTERP163 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV75 : process(INTERP166)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP166);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP165 <= val after tpd_hl;
            when '1' =>
                INTERP165 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV76 : process(INTERP168)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP168);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP167 <= val after tpd_hl;
            when '1' =>
                INTERP167 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV77 : process(INTERP170)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP170);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP169 <= val after tpd_hl;
            when '1' =>
                INTERP169 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV78 : process(INTERP172)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP172);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP171 <= val after tpd_hl;
            when '1' =>
                INTERP171 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV79 : process(INTERP174)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP174);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP173 <= val after tpd_hl;
            when '1' =>
                INTERP173 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV80 : process(INTERP176)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP176);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP175 <= val after tpd_hl;
            when '1' =>
                INTERP175 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV81 : process(INTERP98)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP98);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP177 <= val after tpd_hl;
            when '1' =>
                INTERP177 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV82 : process(INTERP179)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP179);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP178 <= val after tpd_hl;
            when '1' =>
                INTERP178 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV83 : process(INTERP181)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP181);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP180 <= val after tpd_hl;
            when '1' =>
                INTERP180 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV84 : process(INTERP183)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP183);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP182 <= val after tpd_hl;
            when '1' =>
                INTERP182 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV85 : process(INTERP185)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP185);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP184 <= val after tpd_hl;
            when '1' =>
                INTERP184 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV86 : process(INTERP187)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP187);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP186 <= val after tpd_hl;
            when '1' =>
                INTERP186 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV87 : process(INTERP189)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP189);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP188 <= val after tpd_hl;
            when '1' =>
                INTERP188 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV88 : process(INTERP191)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP191);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP190 <= val after tpd_hl;
            when '1' =>
                INTERP190 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV89 : process(INTERP193)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP193);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP192 <= val after tpd_hl;
            when '1' =>
                INTERP192 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV90 : process(INTERP195)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP195);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP194 <= val after tpd_hl;
            when '1' =>
                INTERP194 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV91 : process(INTERP197)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP197);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP196 <= val after tpd_hl;
            when '1' =>
                INTERP196 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV92 : process(INTERP199)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP199);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP198 <= val after tpd_hl;
            when '1' =>
                INTERP198 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV93 : process(INTERP201)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP201);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP200 <= val after tpd_hl;
            when '1' =>
                INTERP200 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND20 : process(INTERP203, INTERP101)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP203 and INTERP101);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP202 <= val after tpd_hl;
            when '1' =>
                INTERP202 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND21 : process(INTERP205, INTERP103)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP205 and INTERP103);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP204 <= val after tpd_hl;
            when '1' =>
                INTERP204 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND22 : process(INTERP207, INTERP105)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP207 and INTERP105);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP206 <= val after tpd_hl;
            when '1' =>
                INTERP206 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND23 : process(INTERP209, INTERP107)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP209 and INTERP107);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP208 <= val after tpd_hl;
            when '1' =>
                INTERP208 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND24 : process(INTERP92, INTERP114)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP92 and INTERP114);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP210 <= val after tpd_hl;
            when '1' =>
                INTERP210 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND25 : process(INTERP212, INTERP116)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP212 and INTERP116);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP211 <= val after tpd_hl;
            when '1' =>
                INTERP211 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND26 : process(INTERP214, INTERP171)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP214 and INTERP171);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP213 <= val after tpd_hl;
            when '1' =>
                INTERP213 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND27 : process(INTERP216, INTERP173)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP216 and INTERP173);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP215 <= val after tpd_hl;
            when '1' =>
                INTERP215 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND28 : process(INTERP218, INTERP177)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP218 and INTERP177);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP217 <= val after tpd_hl;
            when '1' =>
                INTERP217 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND29 : process(INTERP98, INTERP178)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP98 and INTERP178);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP219 <= val after tpd_hl;
            when '1' =>
                INTERP219 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND30 : process(INTERP221, INTERP186)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP221 and INTERP186);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP220 <= val after tpd_hl;
            when '1' =>
                INTERP220 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND31 : process(INTERP223, INTERP188)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP223 and INTERP188);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP222 <= val after tpd_hl;
            when '1' =>
                INTERP222 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND32 : process(INTERP225, INTERP192)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP225 and INTERP192);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP224 <= val after tpd_hl;
            when '1' =>
                INTERP224 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND33 : process(INTERP227, INTERP194)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP227 and INTERP194);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP226 <= val after tpd_hl;
            when '1' =>
                INTERP226 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND34 : process(INTERP229, INTERP198)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP229 and INTERP198);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP228 <= val after tpd_hl;
            when '1' =>
                INTERP228 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND35 : process(INTERP231, INTERP200)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP231 and INTERP200);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP230 <= val after tpd_hl;
            when '1' =>
                INTERP230 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV94 : process(INTERP233)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP233);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP232 <= val after tpd_hl;
            when '1' =>
                INTERP232 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV95 : process(INTERP235)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP235);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP234 <= val after tpd_hl;
            when '1' =>
                INTERP234 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND36 : process(INTERP202, INTERP204)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP202 and INTERP204);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP236 <= val after tpd_hl;
            when '1' =>
                INTERP236 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV96 : process(INTERP238)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP238);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP237 <= val after tpd_hl;
            when '1' =>
                INTERP237 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV97 : process(INTERP240)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP240);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP239 <= val after tpd_hl;
            when '1' =>
                INTERP239 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV98 : process(INTERP242)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP242);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP241 <= val after tpd_hl;
            when '1' =>
                INTERP241 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV99 : process(INTERP244)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP244);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP243 <= val after tpd_hl;
            when '1' =>
                INTERP243 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV100 : process(INTERP246)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP246);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP245 <= val after tpd_hl;
            when '1' =>
                INTERP245 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV101 : process(INTERP248)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP248);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP247 <= val after tpd_hl;
            when '1' =>
                INTERP247 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV102 : process(INTERP250)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP250);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP249 <= val after tpd_hl;
            when '1' =>
                INTERP249 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND37 : process(INTERP206, INTERP208)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP206 and INTERP208);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP251 <= val after tpd_hl;
            when '1' =>
                INTERP251 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV103 : process(INTERP253)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP253);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP252 <= val after tpd_hl;
            when '1' =>
                INTERP252 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND38 : process(INTERP255, INTERP109)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP255 and INTERP109);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP254 <= val after tpd_hl;
            when '1' =>
                INTERP254 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV104 : process(INTERP257)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP257);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP256 <= val after tpd_hl;
            when '1' =>
                INTERP256 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND39 : process(INTERP210, INTERP211)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP210 and INTERP211);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP258 <= val after tpd_hl;
            when '1' =>
                INTERP258 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV105 : process(INTERP119)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP119);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP259 <= val after tpd_hl;
            when '1' =>
                INTERP259 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV106 : process(INTERP120)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP120);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP260 <= val after tpd_hl;
            when '1' =>
                INTERP260 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND40 : process(INTERP139, INTERP145)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP139 and INTERP145);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP261 <= val after tpd_hl;
            when '1' =>
                INTERP261 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND41 : process(INTERP142, INTERP145)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP142 and INTERP145);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP262 <= val after tpd_hl;
            when '1' =>
                INTERP262 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV107 : process(INTERP264)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP264);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP263 <= val after tpd_hl;
            when '1' =>
                INTERP263 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND42 : process(INTERP266, INTERP149)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP266 and INTERP149);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP265 <= val after tpd_hl;
            when '1' =>
                INTERP265 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV108 : process(INTERP268)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP268);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP267 <= val after tpd_hl;
            when '1' =>
                INTERP267 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND43 : process(INTERP270, INTERP151)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP270 and INTERP151);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP269 <= val after tpd_hl;
            when '1' =>
                INTERP269 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV109 : process(INTERP272)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP272);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP271 <= val after tpd_hl;
            when '1' =>
                INTERP271 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND44 : process(INTERP274, INTERP153)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP274 and INTERP153);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP273 <= val after tpd_hl;
            when '1' =>
                INTERP273 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV110 : process(INTERP276)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP276);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP275 <= val after tpd_hl;
            when '1' =>
                INTERP275 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND45 : process(INTERP278, INTERP155)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP278 and INTERP155);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP277 <= val after tpd_hl;
            when '1' =>
                INTERP277 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV111 : process(INTERP280)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP280);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP279 <= val after tpd_hl;
            when '1' =>
                INTERP279 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND46 : process(INTERP282, INTERP157)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP282 and INTERP157);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP281 <= val after tpd_hl;
            when '1' =>
                INTERP281 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV112 : process(INTERP284)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP284);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP283 <= val after tpd_hl;
            when '1' =>
                INTERP283 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND47 : process(INTERP286, INTERP159)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP286 and INTERP159);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP285 <= val after tpd_hl;
            when '1' =>
                INTERP285 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV113 : process(INTERP288)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP288);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP287 <= val after tpd_hl;
            when '1' =>
                INTERP287 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV114 : process(INTERP290)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP290);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP289 <= val after tpd_hl;
            when '1' =>
                INTERP289 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV115 : process(INTERP292)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP292);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP291 <= val after tpd_hl;
            when '1' =>
                INTERP291 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV116 : process(INTERP294)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP294);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP293 <= val after tpd_hl;
            when '1' =>
                INTERP293 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND48 : process(INTERP296, INTERP161)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP296 and INTERP161);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP295 <= val after tpd_hl;
            when '1' =>
                INTERP295 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV117 : process(INTERP298)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP298);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP297 <= val after tpd_hl;
            when '1' =>
                INTERP297 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV118 : process(INTERP300)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP300);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP299 <= val after tpd_hl;
            when '1' =>
                INTERP299 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND49 : process(INTERP302, INTERP163)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP302 and INTERP163);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP301 <= val after tpd_hl;
            when '1' =>
                INTERP301 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV119 : process(INTERP304)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP304);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP303 <= val after tpd_hl;
            when '1' =>
                INTERP303 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND50 : process(INTERP306, INTERP165)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP306 and INTERP165);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP305 <= val after tpd_hl;
            when '1' =>
                INTERP305 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV120 : process(INTERP308)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP308);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP307 <= val after tpd_hl;
            when '1' =>
                INTERP307 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV121 : process(INTERP310)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP310);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP309 <= val after tpd_hl;
            when '1' =>
                INTERP309 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND51 : process(INTERP312, INTERP167)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP312 and INTERP167);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP311 <= val after tpd_hl;
            when '1' =>
                INTERP311 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV122 : process(INTERP314)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP314);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP313 <= val after tpd_hl;
            when '1' =>
                INTERP313 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND52 : process(INTERP316, INTERP169)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP316 and INTERP169);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP315 <= val after tpd_hl;
            when '1' =>
                INTERP315 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND53 : process(INTERP213, INTERP215)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP213 and INTERP215);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP317 <= val after tpd_hl;
            when '1' =>
                INTERP317 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND54 : process(INTERP217, INTERP219)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP217 and INTERP219);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP318 <= val after tpd_hl;
            when '1' =>
                INTERP318 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV123 : process(INTERP320)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP320);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP319 <= val after tpd_hl;
            when '1' =>
                INTERP319 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND55 : process(INTERP322, INTERP182)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP322 and INTERP182);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP321 <= val after tpd_hl;
            when '1' =>
                INTERP321 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV124 : process(INTERP324)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP324);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP323 <= val after tpd_hl;
            when '1' =>
                INTERP323 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV125 : process(INTERP326)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP326);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP325 <= val after tpd_hl;
            when '1' =>
                INTERP325 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND56 : process(INTERP328, INTERP184)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP328 and INTERP184);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP327 <= val after tpd_hl;
            when '1' =>
                INTERP327 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND57 : process(INTERP220, INTERP222)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP220 and INTERP222);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP329 <= val after tpd_hl;
            when '1' =>
                INTERP329 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND58 : process(INTERP224, INTERP226)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP224 and INTERP226);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP330 <= val after tpd_hl;
            when '1' =>
                INTERP330 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND59 : process(INTERP228, INTERP230)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP228 and INTERP230);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP331 <= val after tpd_hl;
            when '1' =>
                INTERP331 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV126 : process(INTERP236)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP236);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP332 <= val after tpd_hl;
            when '1' =>
                INTERP332 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND60 : process(INTERP334, INTERP252)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP334 and INTERP252);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP333 <= val after tpd_hl;
            when '1' =>
                INTERP333 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND61 : process(INTERP336, INTERP263)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP336 and INTERP263);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP335 <= val after tpd_hl;
            when '1' =>
                INTERP335 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND62 : process(INTERP338, INTERP267)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP338 and INTERP267);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP337 <= val after tpd_hl;
            when '1' =>
                INTERP337 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND63 : process(INTERP340, INTERP271)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP340 and INTERP271);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP339 <= val after tpd_hl;
            when '1' =>
                INTERP339 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND64 : process(INTERP342, INTERP275)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP342 and INTERP275);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP341 <= val after tpd_hl;
            when '1' =>
                INTERP341 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND65 : process(INTERP344, INTERP279)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP344 and INTERP279);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP343 <= val after tpd_hl;
            when '1' =>
                INTERP343 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND66 : process(INTERP346, INTERP283)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP346 and INTERP283);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP345 <= val after tpd_hl;
            when '1' =>
                INTERP345 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND67 : process(INTERP348, INTERP293)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP348 and INTERP293);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP347 <= val after tpd_hl;
            when '1' =>
                INTERP347 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND68 : process(INTERP350, INTERP299)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP350 and INTERP299);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP349 <= val after tpd_hl;
            when '1' =>
                INTERP349 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND69 : process(INTERP352, INTERP303)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP352 and INTERP303);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP351 <= val after tpd_hl;
            when '1' =>
                INTERP351 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND70 : process(INTERP354, INTERP309)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP354 and INTERP309);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP353 <= val after tpd_hl;
            when '1' =>
                INTERP353 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV127 : process(INTERP251)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP251);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP355 <= val after tpd_hl;
            when '1' =>
                INTERP355 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND71 : process(INTERP357, INTERP313)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP357 and INTERP313);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP356 <= val after tpd_hl;
            when '1' =>
                INTERP356 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND72 : process(INTERP359, INTERP319)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP359 and INTERP319);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP358 <= val after tpd_hl;
            when '1' =>
                INTERP358 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND73 : process(INTERP361, INTERP325)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP361 and INTERP325);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP360 <= val after tpd_hl;
            when '1' =>
                INTERP360 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV128 : process(INTERP258)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP258);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP362 <= val after tpd_hl;
            when '1' =>
                INTERP362 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND74 : process(INTERP333, INTERP254)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP333 and INTERP254);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP363 <= val after tpd_hl;
            when '1' =>
                INTERP363 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND75 : process(INTERP331, INTERP112)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP331 and INTERP112);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP364 <= val after tpd_hl;
            when '1' =>
                INTERP364 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV129 : process(INTERP331)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP331);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP365 <= val after tpd_hl;
            when '1' =>
                INTERP365 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV130 : process(INTERP367)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP367);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP366 <= val after tpd_hl;
            when '1' =>
                INTERP366 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV131 : process(INTERP369)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP369);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP368 <= val after tpd_hl;
            when '1' =>
                INTERP368 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV132 : process(INTERP371)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP371);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP370 <= val after tpd_hl;
            when '1' =>
                INTERP370 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV133 : process(INTERP373)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP373);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP372 <= val after tpd_hl;
            when '1' =>
                INTERP372 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND76 : process(INTERP335, INTERP265)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP335 and INTERP265);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP374 <= val after tpd_hl;
            when '1' =>
                INTERP374 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND77 : process(INTERP337, INTERP269)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP337 and INTERP269);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP375 <= val after tpd_hl;
            when '1' =>
                INTERP375 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND78 : process(INTERP339, INTERP273)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP339 and INTERP273);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP376 <= val after tpd_hl;
            when '1' =>
                INTERP376 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND79 : process(INTERP341, INTERP277)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP341 and INTERP277);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP377 <= val after tpd_hl;
            when '1' =>
                INTERP377 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND80 : process(INTERP343, INTERP281)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP343 and INTERP281);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP378 <= val after tpd_hl;
            when '1' =>
                INTERP378 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND81 : process(INTERP345, INTERP285)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP345 and INTERP285);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP379 <= val after tpd_hl;
            when '1' =>
                INTERP379 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND82 : process(INTERP347, INTERP295)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP347 and INTERP295);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP380 <= val after tpd_hl;
            when '1' =>
                INTERP380 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND83 : process(INTERP349, INTERP301)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP349 and INTERP301);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP381 <= val after tpd_hl;
            when '1' =>
                INTERP381 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND84 : process(INTERP351, INTERP305)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP351 and INTERP305);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP382 <= val after tpd_hl;
            when '1' =>
                INTERP382 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND85 : process(INTERP353, INTERP311)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP353 and INTERP311);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP383 <= val after tpd_hl;
            when '1' =>
                INTERP383 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND86 : process(INTERP356, INTERP315)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP356 and INTERP315);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP384 <= val after tpd_hl;
            when '1' =>
                INTERP384 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV134 : process(INTERP317)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP317);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP385 <= val after tpd_hl;
            when '1' =>
                INTERP385 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND87 : process(INTERP317, INTERP175)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP317 and INTERP175);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP386 <= val after tpd_hl;
            when '1' =>
                INTERP386 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV135 : process(INTERP318)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP318);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP387 <= val after tpd_hl;
            when '1' =>
                INTERP387 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND88 : process(INTERP318, INTERP180)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP318 and INTERP180);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP388 <= val after tpd_hl;
            when '1' =>
                INTERP388 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND89 : process(INTERP358, INTERP321)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP358 and INTERP321);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP389 <= val after tpd_hl;
            when '1' =>
                INTERP389 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND90 : process(INTERP360, INTERP327)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP360 and INTERP327);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP390 <= val after tpd_hl;
            when '1' =>
                INTERP390 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV136 : process(INTERP329)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP329);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP391 <= val after tpd_hl;
            when '1' =>
                INTERP391 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND91 : process(INTERP329, INTERP190)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP329 and INTERP190);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP392 <= val after tpd_hl;
            when '1' =>
                INTERP392 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV137 : process(INTERP330)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP330);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP393 <= val after tpd_hl;
            when '1' =>
                INTERP393 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND92 : process(INTERP330, INTERP196)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP330 and INTERP196);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP394 <= val after tpd_hl;
            when '1' =>
                INTERP394 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV138 : process(INTERP355)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP355);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP395 <= val after tpd_hl;
            when '1' =>
                INTERP395 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND93 : process(INTERP397, INTERP365)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP397 and INTERP365);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP396 <= val after tpd_hl;
            when '1' =>
                INTERP396 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV139 : process(INTERP362)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP362);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP398 <= val after tpd_hl;
            when '1' =>
                INTERP398 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND94 : process(INTERP400, INTERP385)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP400 and INTERP385);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP399 <= val after tpd_hl;
            when '1' =>
                INTERP399 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND95 : process(INTERP402, INTERP387)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP402 and INTERP387);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP401 <= val after tpd_hl;
            when '1' =>
                INTERP401 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND96 : process(INTERP404, INTERP391)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP404 and INTERP391);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP403 <= val after tpd_hl;
            when '1' =>
                INTERP403 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND97 : process(INTERP406, INTERP393)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP406 and INTERP393);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP405 <= val after tpd_hl;
            when '1' =>
                INTERP405 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV140 : process(INTERP363)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP363);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP407 <= val after tpd_hl;
            when '1' =>
                INTERP407 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND98 : process(INTERP375, INTERP232)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP375 and INTERP232);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP408 <= val after tpd_hl;
            when '1' =>
                INTERP408 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV141 : process(INTERP375)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP375);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP409 <= val after tpd_hl;
            when '1' =>
                INTERP409 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND99 : process(INTERP374, INTERP234)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP374 and INTERP234);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP410 <= val after tpd_hl;
            when '1' =>
                INTERP410 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV142 : process(INTERP374)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP374);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP411 <= val after tpd_hl;
            when '1' =>
                INTERP411 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND100 : process(INTERP376, INTERP237)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP376 and INTERP237);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP412 <= val after tpd_hl;
            when '1' =>
                INTERP412 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV143 : process(INTERP376)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP376);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP413 <= val after tpd_hl;
            when '1' =>
                INTERP413 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND101 : process(INTERP377, INTERP239)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP377 and INTERP239);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP414 <= val after tpd_hl;
            when '1' =>
                INTERP414 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV144 : process(INTERP377)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP377);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP415 <= val after tpd_hl;
            when '1' =>
                INTERP415 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND102 : process(INTERP379, INTERP241)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP379 and INTERP241);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP416 <= val after tpd_hl;
            when '1' =>
                INTERP416 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV145 : process(INTERP379)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP379);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP417 <= val after tpd_hl;
            when '1' =>
                INTERP417 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND103 : process(INTERP378, INTERP243)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP378 and INTERP243);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP418 <= val after tpd_hl;
            when '1' =>
                INTERP418 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV146 : process(INTERP378)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP378);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP419 <= val after tpd_hl;
            when '1' =>
                INTERP419 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND104 : process(INTERP381, INTERP247)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP381 and INTERP247);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP420 <= val after tpd_hl;
            when '1' =>
                INTERP420 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV147 : process(INTERP381)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP381);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP421 <= val after tpd_hl;
            when '1' =>
                INTERP421 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND105 : process(INTERP383, INTERP249)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP383 and INTERP249);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP422 <= val after tpd_hl;
            when '1' =>
                INTERP422 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV148 : process(INTERP383)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP383);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP423 <= val after tpd_hl;
            when '1' =>
                INTERP423 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV149 : process(INTERP384)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP384);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP424 <= val after tpd_hl;
            when '1' =>
                INTERP424 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND106 : process(INTERP390, INTERP256)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP390 and INTERP256);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP425 <= val after tpd_hl;
            when '1' =>
                INTERP425 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV150 : process(INTERP390)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP390);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP426 <= val after tpd_hl;
            when '1' =>
                INTERP426 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND107 : process(INTERP364, INTERP396)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP364 and INTERP396);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP427 <= val after tpd_hl;
            when '1' =>
                INTERP427 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV151 : process(INTERP380)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP380);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP428 <= val after tpd_hl;
            when '1' =>
                INTERP428 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND108 : process(INTERP380, INTERP297)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP380 and INTERP297);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP429 <= val after tpd_hl;
            when '1' =>
                INTERP429 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV152 : process(INTERP382)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP382);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP430 <= val after tpd_hl;
            when '1' =>
                INTERP430 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND109 : process(INTERP382, INTERP307)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP382 and INTERP307);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP431 <= val after tpd_hl;
            when '1' =>
                INTERP431 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND110 : process(INTERP386, INTERP399)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP386 and INTERP399);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP432 <= val after tpd_hl;
            when '1' =>
                INTERP432 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV153 : process(INTERP389)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP389);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP433 <= val after tpd_hl;
            when '1' =>
                INTERP433 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND111 : process(INTERP389, INTERP323)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP389 and INTERP323);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP434 <= val after tpd_hl;
            when '1' =>
                INTERP434 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND112 : process(INTERP388, INTERP401)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP388 and INTERP401);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP435 <= val after tpd_hl;
            when '1' =>
                INTERP435 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND113 : process(INTERP394, INTERP405)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP394 and INTERP405);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP436 <= val after tpd_hl;
            when '1' =>
                INTERP436 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND114 : process(INTERP392, INTERP403)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP392 and INTERP403);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP437 <= val after tpd_hl;
            when '1' =>
                INTERP437 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND115 : process(INTERP439, INTERP409)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP439 and INTERP409);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP438 <= val after tpd_hl;
            when '1' =>
                INTERP438 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND116 : process(INTERP441, INTERP411)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP441 and INTERP411);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP440 <= val after tpd_hl;
            when '1' =>
                INTERP440 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND117 : process(INTERP443, INTERP413)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP443 and INTERP413);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP442 <= val after tpd_hl;
            when '1' =>
                INTERP442 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV154 : process(INTERP445)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP445);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP444 <= val after tpd_hl;
            when '1' =>
                INTERP444 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV155 : process(INTERP447)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP447);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP446 <= val after tpd_hl;
            when '1' =>
                INTERP446 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND118 : process(INTERP449, INTERP415)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP449 and INTERP415);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP448 <= val after tpd_hl;
            when '1' =>
                INTERP448 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND119 : process(INTERP451, INTERP417)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP451 and INTERP417);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP450 <= val after tpd_hl;
            when '1' =>
                INTERP450 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND120 : process(INTERP453, INTERP419)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP453 and INTERP419);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP452 <= val after tpd_hl;
            when '1' =>
                INTERP452 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND121 : process(INTERP455, INTERP421)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP455 and INTERP421);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP454 <= val after tpd_hl;
            when '1' =>
                INTERP454 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND122 : process(INTERP457, INTERP423)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP457 and INTERP423);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP456 <= val after tpd_hl;
            when '1' =>
                INTERP456 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND123 : process(INTERP459, INTERP426)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP459 and INTERP426);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP458 <= val after tpd_hl;
            when '1' =>
                INTERP458 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV156 : process(INTERP407)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP407);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP460 <= val after tpd_hl;
            when '1' =>
                INTERP460 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND124 : process(INTERP462, INTERP428)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP462 and INTERP428);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP461 <= val after tpd_hl;
            when '1' =>
                INTERP461 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND125 : process(INTERP464, INTERP430)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP464 and INTERP430);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP463 <= val after tpd_hl;
            when '1' =>
                INTERP463 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND126 : process(INTERP466, INTERP433)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP466 and INTERP433);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP465 <= val after tpd_hl;
            when '1' =>
                INTERP465 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV157 : process(INTERP427)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP427);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP467 <= val after tpd_hl;
            when '1' =>
                INTERP467 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND127 : process(INTERP408, INTERP438)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP408 and INTERP438);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP468 <= val after tpd_hl;
            when '1' =>
                INTERP468 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND128 : process(INTERP410, INTERP440)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP410 and INTERP440);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP469 <= val after tpd_hl;
            when '1' =>
                INTERP469 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND129 : process(INTERP412, INTERP442)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP412 and INTERP442);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP470 <= val after tpd_hl;
            when '1' =>
                INTERP470 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND130 : process(INTERP414, INTERP448)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP414 and INTERP448);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP471 <= val after tpd_hl;
            when '1' =>
                INTERP471 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND131 : process(INTERP416, INTERP450)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP416 and INTERP450);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP472 <= val after tpd_hl;
            when '1' =>
                INTERP472 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND132 : process(INTERP418, INTERP452)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP418 and INTERP452);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP473 <= val after tpd_hl;
            when '1' =>
                INTERP473 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND133 : process(INTERP420, INTERP454)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP420 and INTERP454);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP474 <= val after tpd_hl;
            when '1' =>
                INTERP474 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND134 : process(INTERP422, INTERP456)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP422 and INTERP456);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP475 <= val after tpd_hl;
            when '1' =>
                INTERP475 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV158 : process(INTERP432)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP432);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP476 <= val after tpd_hl;
            when '1' =>
                INTERP476 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND135 : process(INTERP425, INTERP458)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP425 and INTERP458);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP477 <= val after tpd_hl;
            when '1' =>
                INTERP477 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV159 : process(INTERP435)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP435);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP478 <= val after tpd_hl;
            when '1' =>
                INTERP478 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV160 : process(INTERP436)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP436);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP479 <= val after tpd_hl;
            when '1' =>
                INTERP479 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV161 : process(INTERP437)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP437);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP480 <= val after tpd_hl;
            when '1' =>
                INTERP480 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND136 : process(INTERP431, INTERP463)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP431 and INTERP463);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP481 <= val after tpd_hl;
            when '1' =>
                INTERP481 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND137 : process(INTERP429, INTERP461)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP429 and INTERP461);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP482 <= val after tpd_hl;
            when '1' =>
                INTERP482 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND138 : process(INTERP434, INTERP465)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP434 and INTERP465);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP483 <= val after tpd_hl;
            when '1' =>
                INTERP483 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV162 : process(INTERP468)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP468);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP484 <= val after tpd_hl;
            when '1' =>
                INTERP484 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV163 : process(INTERP472)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP472);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP485 <= val after tpd_hl;
            when '1' =>
                INTERP485 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV164 : process(INTERP474)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP474);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP486 <= val after tpd_hl;
            when '1' =>
                INTERP486 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV165 : process(INTERP471)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP471);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP487 <= val after tpd_hl;
            when '1' =>
                INTERP487 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND139 : process(INTERP437, INTERP479)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP437 and INTERP479);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP488 <= val after tpd_hl;
            when '1' =>
                INTERP488 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND140 : process(INTERP436, INTERP480)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP436 and INTERP480);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP489 <= val after tpd_hl;
            when '1' =>
                INTERP489 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV166 : process(INTERP467)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP467);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP490 <= val after tpd_hl;
            when '1' =>
                INTERP490 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV167 : process(INTERP475)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP475);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP491 <= val after tpd_hl;
            when '1' =>
                INTERP491 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV168 : process(INTERP477)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP477);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP492 <= val after tpd_hl;
            when '1' =>
                INTERP492 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV169 : process(INTERP481)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP481);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP493 <= val after tpd_hl;
            when '1' =>
                INTERP493 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV170 : process(INTERP482)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP482);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP494 <= val after tpd_hl;
            when '1' =>
                INTERP494 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND141 : process(INTERP483, INTERP478)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP483 and INTERP478);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP495 <= val after tpd_hl;
            when '1' =>
                INTERP495 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV171 : process(INTERP483)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP483);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP496 <= val after tpd_hl;
            when '1' =>
                INTERP496 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND142 : process(INTERP488, INTERP489)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP488 and INTERP489);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP497 <= val after tpd_hl;
            when '1' =>
                INTERP497 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV172 : process(INTERP491)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP491);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP498 <= val after tpd_hl;
            when '1' =>
                INTERP498 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND143 : process(INTERP435, INTERP496)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP435 and INTERP496);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP499 <= val after tpd_hl;
            when '1' =>
                INTERP499 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND144 : process(INTERP492, INTERP490)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP492 and INTERP490);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP500 <= val after tpd_hl;
            when '1' =>
                INTERP500 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV173 : process(INTERP492)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP492);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP501 <= val after tpd_hl;
            when '1' =>
                INTERP501 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND145 : process(INTERP497, INTERP111)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP497 and INTERP111);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP502 <= val after tpd_hl;
            when '1' =>
                INTERP502 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV174 : process(INTERP497)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP497);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP503 <= val after tpd_hl;
            when '1' =>
                INTERP503 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV175 : process(INTERP505)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP505);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP504 <= val after tpd_hl;
            when '1' =>
                INTERP504 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV176 : process(INTERP507)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP507);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP506 <= val after tpd_hl;
            when '1' =>
                INTERP506 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND146 : process(INTERP509, INTERP287)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP509 and INTERP287);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP508 <= val after tpd_hl;
            when '1' =>
                INTERP508 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV177 : process(INTERP511)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP511);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP510 <= val after tpd_hl;
            when '1' =>
                INTERP510 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND147 : process(INTERP513, INTERP291)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP513 and INTERP291);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP512 <= val after tpd_hl;
            when '1' =>
                INTERP512 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV178 : process(INTERP515)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP515);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP514 <= val after tpd_hl;
            when '1' =>
                INTERP514 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV179 : process(INTERP517)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP517);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP516 <= val after tpd_hl;
            when '1' =>
                INTERP516 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV180 : process(INTERP519)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP519);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP518 <= val after tpd_hl;
            when '1' =>
                INTERP518 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND148 : process(INTERP495, INTERP499)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP495 and INTERP499);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP520 <= val after tpd_hl;
            when '1' =>
                INTERP520 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND149 : process(INTERP467, INTERP501)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP467 and INTERP501);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP521 <= val after tpd_hl;
            when '1' =>
                INTERP521 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND150 : process(INTERP90, INTERP503)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP90 and INTERP503);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP522 <= val after tpd_hl;
            when '1' =>
                INTERP522 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV181 : process(INTERP524)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP524);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP523 <= val after tpd_hl;
            when '1' =>
                INTERP523 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND151 : process(INTERP526, INTERP504)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP526 and INTERP504);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP525 <= val after tpd_hl;
            when '1' =>
                INTERP525 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV182 : process(INTERP528)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP528);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP527 <= val after tpd_hl;
            when '1' =>
                INTERP527 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND152 : process(INTERP530, INTERP506)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP530 and INTERP506);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP529 <= val after tpd_hl;
            when '1' =>
                INTERP529 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV183 : process(INTERP532)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP532);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP531 <= val after tpd_hl;
            when '1' =>
                INTERP531 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND153 : process(INTERP534, INTERP510)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP534 and INTERP510);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP533 <= val after tpd_hl;
            when '1' =>
                INTERP533 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND154 : process(INTERP536, INTERP514)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP536 and INTERP514);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP535 <= val after tpd_hl;
            when '1' =>
                INTERP535 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND155 : process(INTERP538, INTERP494)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP538 and INTERP494);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP537 <= val after tpd_hl;
            when '1' =>
                INTERP537 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV184 : process(INTERP540)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP540);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP539 <= val after tpd_hl;
            when '1' =>
                INTERP539 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND156 : process(INTERP500, INTERP521)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP500 and INTERP521);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP541 <= val after tpd_hl;
            when '1' =>
                INTERP541 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV185 : process(INTERP543)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP543);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP542 <= val after tpd_hl;
            when '1' =>
                INTERP542 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV186 : process(INTERP545)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP545);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP544 <= val after tpd_hl;
            when '1' =>
                INTERP544 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV187 : process(INTERP547)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP547);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP546 <= val after tpd_hl;
            when '1' =>
                INTERP546 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND157 : process(INTERP520, INTERP476)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP520 and INTERP476);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP548 <= val after tpd_hl;
            when '1' =>
                INTERP548 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV188 : process(INTERP520)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP520);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP549 <= val after tpd_hl;
            when '1' =>
                INTERP549 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND158 : process(INTERP502, INTERP522)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP502 and INTERP522);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP550 <= val after tpd_hl;
            when '1' =>
                INTERP550 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND159 : process(INTERP552, INTERP527)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP552 and INTERP527);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP551 <= val after tpd_hl;
            when '1' =>
                INTERP551 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND160 : process(INTERP554, INTERP531)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP554 and INTERP531);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP553 <= val after tpd_hl;
            when '1' =>
                INTERP553 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND161 : process(INTERP508, INTERP533)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP508 and INTERP533);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP555 <= val after tpd_hl;
            when '1' =>
                INTERP555 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND162 : process(INTERP512, INTERP535)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP512 and INTERP535);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP556 <= val after tpd_hl;
            when '1' =>
                INTERP556 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND163 : process(INTERP482, INTERP539)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP482 and INTERP539);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP557 <= val after tpd_hl;
            when '1' =>
                INTERP557 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV189 : process(INTERP559)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP559);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP558 <= val after tpd_hl;
            when '1' =>
                INTERP558 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND164 : process(INTERP561, INTERP542)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP561 and INTERP542);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP560 <= val after tpd_hl;
            when '1' =>
                INTERP560 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV190 : process(INTERP563)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP563);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP562 <= val after tpd_hl;
            when '1' =>
                INTERP562 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND165 : process(INTERP565, INTERP546)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP565 and INTERP546);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP564 <= val after tpd_hl;
            when '1' =>
                INTERP564 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV191 : process(INTERP567)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP567);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP566 <= val after tpd_hl;
            when '1' =>
                INTERP566 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND166 : process(INTERP432, INTERP549)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP432 and INTERP549);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP568 <= val after tpd_hl;
            when '1' =>
                INTERP568 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND167 : process(INTERP541, INTERP398)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP541 and INTERP398);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP569 <= val after tpd_hl;
            when '1' =>
                INTERP569 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV192 : process(INTERP541)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP541);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP570 <= val after tpd_hl;
            when '1' =>
                INTERP570 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND168 : process(INTERP525, INTERP551)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP525 and INTERP551);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP571 <= val after tpd_hl;
            when '1' =>
                INTERP571 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND169 : process(INTERP529, INTERP553)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP529 and INTERP553);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP572 <= val after tpd_hl;
            when '1' =>
                INTERP572 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV193 : process(INTERP574)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP574);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP573 <= val after tpd_hl;
            when '1' =>
                INTERP573 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND170 : process(INTERP576, INTERP516)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP576 and INTERP516);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP575 <= val after tpd_hl;
            when '1' =>
                INTERP575 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV194 : process(INTERP578)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP578);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP577 <= val after tpd_hl;
            when '1' =>
                INTERP577 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV195 : process(INTERP580)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP580);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP579 <= val after tpd_hl;
            when '1' =>
                INTERP579 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND171 : process(INTERP582, INTERP518)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP582 and INTERP518);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP581 <= val after tpd_hl;
            when '1' =>
                INTERP581 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND172 : process(INTERP537, INTERP557)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP537 and INTERP557);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP583 <= val after tpd_hl;
            when '1' =>
                INTERP583 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND173 : process(INTERP585, INTERP558)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP585 and INTERP558);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP584 <= val after tpd_hl;
            when '1' =>
                INTERP584 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND174 : process(INTERP587, INTERP562)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP587 and INTERP562);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP586 <= val after tpd_hl;
            when '1' =>
                INTERP586 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND175 : process(INTERP556, INTERP245)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP556 and INTERP245);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP588 <= val after tpd_hl;
            when '1' =>
                INTERP588 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV196 : process(INTERP556)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP556);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP589 <= val after tpd_hl;
            when '1' =>
                INTERP589 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND176 : process(INTERP548, INTERP568)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP548 and INTERP568);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP590 <= val after tpd_hl;
            when '1' =>
                INTERP590 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND177 : process(INTERP362, INTERP570)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP362 and INTERP570);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP591 <= val after tpd_hl;
            when '1' =>
                INTERP591 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND178 : process(INTERP550, INTERP28)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP550 and INTERP28);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP592 <= val after tpd_hl;
            when '1' =>
                INTERP592 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV197 : process(INTERP555)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP555);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP593 <= val after tpd_hl;
            when '1' =>
                INTERP593 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND179 : process(INTERP555, INTERP289)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP555 and INTERP289);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP594 <= val after tpd_hl;
            when '1' =>
                INTERP594 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND180 : process(INTERP596, INTERP573)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP596 and INTERP573);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP595 <= val after tpd_hl;
            when '1' =>
                INTERP595 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND181 : process(INTERP598, INTERP579)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP598 and INTERP579);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP597 <= val after tpd_hl;
            when '1' =>
                INTERP597 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND182 : process(INTERP584, INTERP560)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP584 and INTERP560);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP599 <= val after tpd_hl;
            when '1' =>
                INTERP599 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND183 : process(INTERP586, INTERP564)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP586 and INTERP564);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP600 <= val after tpd_hl;
            when '1' =>
                INTERP600 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND184 : process(INTERP572, INTERP444)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP572 and INTERP444);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP601 <= val after tpd_hl;
            when '1' =>
                INTERP601 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV198 : process(INTERP572)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP572);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP602 <= val after tpd_hl;
            when '1' =>
                INTERP602 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND185 : process(INTERP571, INTERP446)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP571 and INTERP446);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP603 <= val after tpd_hl;
            when '1' =>
                INTERP603 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV199 : process(INTERP571)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP571);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP604 <= val after tpd_hl;
            when '1' =>
                INTERP604 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND186 : process(INTERP606, INTERP589)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP606 and INTERP589);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP605 <= val after tpd_hl;
            when '1' =>
                INTERP605 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND187 : process(INTERP583, INTERP395)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP583 and INTERP395);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP607 <= val after tpd_hl;
            when '1' =>
                INTERP607 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV200 : process(INTERP583)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP583);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP608 <= val after tpd_hl;
            when '1' =>
                INTERP608 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND188 : process(INTERP569, INTERP591)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP569 and INTERP591);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP609 <= val after tpd_hl;
            when '1' =>
                INTERP609 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND189 : process(INTERP611, INTERP593)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP611 and INTERP593);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP610 <= val after tpd_hl;
            when '1' =>
                INTERP610 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND190 : process(INTERP595, INTERP575)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP595 and INTERP575);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP612 <= val after tpd_hl;
            when '1' =>
                INTERP612 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND191 : process(INTERP597, INTERP581)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP597 and INTERP581);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP613 <= val after tpd_hl;
            when '1' =>
                INTERP613 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND192 : process(INTERP615, INTERP602)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP615 and INTERP602);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP614 <= val after tpd_hl;
            when '1' =>
                INTERP614 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND193 : process(INTERP617, INTERP604)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP617 and INTERP604);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP616 <= val after tpd_hl;
            when '1' =>
                INTERP616 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND194 : process(INTERP588, INTERP605)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP588 and INTERP605);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP618 <= val after tpd_hl;
            when '1' =>
                INTERP618 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND195 : process(INTERP355, INTERP608)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP355 and INTERP608);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP619 <= val after tpd_hl;
            when '1' =>
                INTERP619 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND196 : process(INTERP600, INTERP523)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP600 and INTERP523);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP620 <= val after tpd_hl;
            when '1' =>
                INTERP620 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV201 : process(INTERP600)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP600);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP621 <= val after tpd_hl;
            when '1' =>
                INTERP621 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV202 : process(INTERP623)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP623);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP622 <= val after tpd_hl;
            when '1' =>
                INTERP622 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND197 : process(INTERP590, INTERP28)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP590 and INTERP28);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP624 <= val after tpd_hl;
            when '1' =>
                INTERP624 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV203 : process(INTERP599)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP599);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP625 <= val after tpd_hl;
            when '1' =>
                INTERP625 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND198 : process(INTERP599, INTERP544)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP599 and INTERP544);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP626 <= val after tpd_hl;
            when '1' =>
                INTERP626 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND199 : process(INTERP594, INTERP610)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP594 and INTERP610);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP627 <= val after tpd_hl;
            when '1' =>
                INTERP627 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND200 : process(INTERP601, INTERP614)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP601 and INTERP614);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP628 <= val after tpd_hl;
            when '1' =>
                INTERP628 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND201 : process(INTERP603, INTERP616)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP603 and INTERP616);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP629 <= val after tpd_hl;
            when '1' =>
                INTERP629 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND202 : process(INTERP613, INTERP566)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP613 and INTERP566);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP630 <= val after tpd_hl;
            when '1' =>
                INTERP630 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV204 : process(INTERP613)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP613);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP631 <= val after tpd_hl;
            when '1' =>
                INTERP631 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND203 : process(INTERP607, INTERP619)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP607 and INTERP619);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP632 <= val after tpd_hl;
            when '1' =>
                INTERP632 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND204 : process(INTERP634, INTERP621)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP634 and INTERP621);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP633 <= val after tpd_hl;
            when '1' =>
                INTERP633 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND205 : process(INTERP609, INTERP28)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP609 and INTERP28);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP635 <= val after tpd_hl;
            when '1' =>
                INTERP635 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV205 : process(INTERP612)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP612);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP636 <= val after tpd_hl;
            when '1' =>
                INTERP636 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND206 : process(INTERP612, INTERP577)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP612 and INTERP577);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP637 <= val after tpd_hl;
            when '1' =>
                INTERP637 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND207 : process(INTERP639, INTERP625)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP639 and INTERP625);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP638 <= val after tpd_hl;
            when '1' =>
                INTERP638 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV206 : process(INTERP618)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP618);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP640 <= val after tpd_hl;
            when '1' =>
                INTERP640 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV207 : process(INTERP628)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP628);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP641 <= val after tpd_hl;
            when '1' =>
                INTERP641 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND208 : process(INTERP643, INTERP631)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP643 and INTERP631);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP642 <= val after tpd_hl;
            when '1' =>
                INTERP642 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV208 : process(INTERP632)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP632);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP644 <= val after tpd_hl;
            when '1' =>
                INTERP644 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND209 : process(INTERP620, INTERP633)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP620 and INTERP633);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP645 <= val after tpd_hl;
            when '1' =>
                INTERP645 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV209 : process(INTERP647)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP647);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP646 <= val after tpd_hl;
            when '1' =>
                INTERP646 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND210 : process(INTERP649, INTERP135)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP649 and INTERP135);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP648 <= val after tpd_hl;
            when '1' =>
                INTERP648 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV210 : process(INTERP651)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP651);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP650 <= val after tpd_hl;
            when '1' =>
                INTERP650 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND211 : process(INTERP653, INTERP137)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP653 and INTERP137);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP652 <= val after tpd_hl;
            when '1' =>
                INTERP652 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV211 : process(INTERP655)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP655);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP654 <= val after tpd_hl;
            when '1' =>
                INTERP654 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV212 : process(INTERP627)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP627);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP656 <= val after tpd_hl;
            when '1' =>
                INTERP656 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND212 : process(INTERP658, INTERP636)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP658 and INTERP636);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP657 <= val after tpd_hl;
            when '1' =>
                INTERP657 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND213 : process(INTERP626, INTERP638)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP626 and INTERP638);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP659 <= val after tpd_hl;
            when '1' =>
                INTERP659 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND214 : process(INTERP630, INTERP642)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP630 and INTERP642);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP660 <= val after tpd_hl;
            when '1' =>
                INTERP660 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV213 : process(INTERP640)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP640);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP661 <= val after tpd_hl;
            when '1' =>
                INTERP661 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV214 : process(INTERP663)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP663);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP662 <= val after tpd_hl;
            when '1' =>
                INTERP662 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND215 : process(INTERP665, INTERP650)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP665 and INTERP650);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP664 <= val after tpd_hl;
            when '1' =>
                INTERP664 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND216 : process(INTERP667, INTERP654)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP667 and INTERP654);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP666 <= val after tpd_hl;
            when '1' =>
                INTERP666 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV215 : process(INTERP645)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP645);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP668 <= val after tpd_hl;
            when '1' =>
                INTERP668 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND217 : process(INTERP637, INTERP657)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP637 and INTERP657);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP669 <= val after tpd_hl;
            when '1' =>
                INTERP669 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND11 : process(INTERP641, INTERP81)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP641 and INTERP81;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP670 <= val after tpd_hl;
            when '1' =>
                INTERP670 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND12 : process(INTERP83, INTERP644)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP83 and INTERP644;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP671 <= val after tpd_hl;
            when '1' =>
                INTERP671 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND218 : process(INTERP673, INTERP131)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP673 and INTERP131);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP672 <= val after tpd_hl;
            when '1' =>
                INTERP672 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV216 : process(INTERP675)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP675);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP674 <= val after tpd_hl;
            when '1' =>
                INTERP674 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND219 : process(INTERP677, INTERP133)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP677 and INTERP133);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP676 <= val after tpd_hl;
            when '1' =>
                INTERP676 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV217 : process(INTERP679)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP679);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP678 <= val after tpd_hl;
            when '1' =>
                INTERP678 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND220 : process(INTERP648, INTERP664)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP648 and INTERP664);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP680 <= val after tpd_hl;
            when '1' =>
                INTERP680 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND221 : process(INTERP652, INTERP666)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP652 and INTERP666);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP681 <= val after tpd_hl;
            when '1' =>
                INTERP681 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV218 : process(INTERP659)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP659);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP682 <= val after tpd_hl;
            when '1' =>
                INTERP682 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV219 : process(INTERP660)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP660);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP683 <= val after tpd_hl;
            when '1' =>
                INTERP683 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV220 : process(INTERP685)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP685);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP684 <= val after tpd_hl;
            when '1' =>
                INTERP684 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND222 : process(INTERP687, INTERP661)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP687 and INTERP661);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP686 <= val after tpd_hl;
            when '1' =>
                INTERP686 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV221 : process(INTERP668)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP668);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP688 <= val after tpd_hl;
            when '1' =>
                INTERP688 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND223 : process(INTERP668, INTERP460)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP668 and INTERP460);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP689 <= val after tpd_hl;
            when '1' =>
                INTERP689 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND224 : process(INTERP691, INTERP370)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP691 and INTERP370);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP690 <= val after tpd_hl;
            when '1' =>
                INTERP690 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV222 : process(INTERP693)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP693);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP692 <= val after tpd_hl;
            when '1' =>
                INTERP692 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND225 : process(INTERP695, INTERP372)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP695 and INTERP372);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP694 <= val after tpd_hl;
            when '1' =>
                INTERP694 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV223 : process(INTERP697)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP697);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP696 <= val after tpd_hl;
            when '1' =>
                INTERP696 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND226 : process(INTERP699, INTERP674)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP699 and INTERP674);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP698 <= val after tpd_hl;
            when '1' =>
                INTERP698 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND227 : process(INTERP701, INTERP678)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP701 and INTERP678);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP700 <= val after tpd_hl;
            when '1' =>
                INTERP700 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV224 : process(INTERP680)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP680);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP702 <= val after tpd_hl;
            when '1' =>
                INTERP702 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV225 : process(INTERP704)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP704);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP703 <= val after tpd_hl;
            when '1' =>
                INTERP703 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND228 : process(INTERP706, INTERP656)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP706 and INTERP656);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP705 <= val after tpd_hl;
            when '1' =>
                INTERP705 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV226 : process(INTERP669)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP669);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP707 <= val after tpd_hl;
            when '1' =>
                INTERP707 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND229 : process(INTERP669, INTERP498)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP669 and INTERP498);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP708 <= val after tpd_hl;
            when '1' =>
                INTERP708 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV227 : process(INTERP670)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP670);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP709 <= val after tpd_hl;
            when '1' =>
                INTERP709 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV228 : process(INTERP671)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP671);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP710 <= val after tpd_hl;
            when '1' =>
                INTERP710 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND230 : process(INTERP640, INTERP684)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP640 and INTERP684);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP711 <= val after tpd_hl;
            when '1' =>
                INTERP711 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV229 : process(INTERP683)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP683);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP712 <= val after tpd_hl;
            when '1' =>
                INTERP712 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND231 : process(INTERP683, INTERP493)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP683 and INTERP493);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP713 <= val after tpd_hl;
            when '1' =>
                INTERP713 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND232 : process(INTERP407, INTERP688)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP407 and INTERP688);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP714 <= val after tpd_hl;
            when '1' =>
                INTERP714 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND233 : process(INTERP716, INTERP692)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP716 and INTERP692);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP715 <= val after tpd_hl;
            when '1' =>
                INTERP715 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND234 : process(INTERP718, INTERP696)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP718 and INTERP696);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP717 <= val after tpd_hl;
            when '1' =>
                INTERP717 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND235 : process(INTERP672, INTERP698)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP672 and INTERP698);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP719 <= val after tpd_hl;
            when '1' =>
                INTERP719 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND236 : process(INTERP676, INTERP700)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP676 and INTERP700);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP720 <= val after tpd_hl;
            when '1' =>
                INTERP720 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV230 : process(INTERP681)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP681);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP721 <= val after tpd_hl;
            when '1' =>
                INTERP721 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND237 : process(INTERP627, INTERP703)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP627 and INTERP703);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP722 <= val after tpd_hl;
            when '1' =>
                INTERP722 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND238 : process(INTERP491, INTERP707)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP491 and INTERP707);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP723 <= val after tpd_hl;
            when '1' =>
                INTERP723 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND239 : process(INTERP711, INTERP686)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP711 and INTERP686);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP724 <= val after tpd_hl;
            when '1' =>
                INTERP724 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND240 : process(INTERP481, INTERP712)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP481 and INTERP712);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP725 <= val after tpd_hl;
            when '1' =>
                INTERP725 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND241 : process(INTERP714, INTERP689)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP714 and INTERP689);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP726 <= val after tpd_hl;
            when '1' =>
                INTERP726 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND242 : process(INTERP690, INTERP715)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP690 and INTERP715);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP727 <= val after tpd_hl;
            when '1' =>
                INTERP727 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND243 : process(INTERP694, INTERP717)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP694 and INTERP717);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP728 <= val after tpd_hl;
            when '1' =>
                INTERP728 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV231 : process(INTERP719)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP719);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP729 <= val after tpd_hl;
            when '1' =>
                INTERP729 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND244 : process(INTERP722, INTERP705)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP722 and INTERP705);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP730 <= val after tpd_hl;
            when '1' =>
                INTERP730 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND245 : process(INTERP723, INTERP708)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP723 and INTERP708);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP731 <= val after tpd_hl;
            when '1' =>
                INTERP731 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV232 : process(INTERP724)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP724);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP732 <= val after tpd_hl;
            when '1' =>
                INTERP732 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND246 : process(INTERP725, INTERP713)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP725 and INTERP713);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP733 <= val after tpd_hl;
            when '1' =>
                INTERP733 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND247 : process(INTERP726, INTERP28)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP726 and INTERP28);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP734 <= val after tpd_hl;
            when '1' =>
                INTERP734 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV233 : process(INTERP727)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP727);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP735 <= val after tpd_hl;
            when '1' =>
                INTERP735 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV234 : process(INTERP720)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP720);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP736 <= val after tpd_hl;
            when '1' =>
                INTERP736 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV235 : process(INTERP730)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP730);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP737 <= val after tpd_hl;
            when '1' =>
                INTERP737 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV236 : process(INTERP731)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP731);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP738 <= val after tpd_hl;
            when '1' =>
                INTERP738 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND248 : process(INTERP732, INTERP28)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP732 and INTERP28);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP739 <= val after tpd_hl;
            when '1' =>
                INTERP739 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND249 : process(INTERP733, INTERP28)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP733 and INTERP28);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP740 <= val after tpd_hl;
            when '1' =>
                INTERP740 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV237 : process(INTERP728)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP728);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP741 <= val after tpd_hl;
            when '1' =>
                INTERP741 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND13 : process(INTERP721, INTERP736)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP721 and INTERP736;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP742 <= val after tpd_hl;
            when '1' =>
                INTERP742 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND14 : process(INTERP744, INTERP736)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP744 and INTERP736;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP743 <= val after tpd_hl;
            when '1' =>
                INTERP743 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND15 : process(INTERP721, INTERP746)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP721 and INTERP746;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP745 <= val after tpd_hl;
            when '1' =>
                INTERP745 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND16 : process(INTERP748, INTERP749)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP748 and INTERP749;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP747 <= val after tpd_hl;
            when '1' =>
                INTERP747 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND250 : process(INTERP751, INTERP127)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP751 and INTERP127);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP750 <= val after tpd_hl;
            when '1' =>
                INTERP750 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV238 : process(INTERP753)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP753);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP752 <= val after tpd_hl;
            when '1' =>
                INTERP752 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND251 : process(INTERP755, INTERP129)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP755 and INTERP129);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP754 <= val after tpd_hl;
            when '1' =>
                INTERP754 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV239 : process(INTERP757)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP757);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP756 <= val after tpd_hl;
            when '1' =>
                INTERP756 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND252 : process(INTERP759, INTERP366)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP759 and INTERP366);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP758 <= val after tpd_hl;
            when '1' =>
                INTERP758 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV240 : process(INTERP761)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP761);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP760 <= val after tpd_hl;
            when '1' =>
                INTERP760 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND253 : process(INTERP763, INTERP368)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP763 and INTERP368);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP762 <= val after tpd_hl;
            when '1' =>
                INTERP762 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV241 : process(INTERP765)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP765);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP764 <= val after tpd_hl;
            when '1' =>
                INTERP764 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND254 : process(INTERP767, INTERP123)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP767 and INTERP123);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP766 <= val after tpd_hl;
            when '1' =>
                INTERP766 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV242 : process(INTERP769)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP769);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP768 <= val after tpd_hl;
            when '1' =>
                INTERP768 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND255 : process(INTERP771, INTERP125)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP771 and INTERP125);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP770 <= val after tpd_hl;
            when '1' =>
                INTERP770 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV243 : process(INTERP773)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP773);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP772 <= val after tpd_hl;
            when '1' =>
                INTERP772 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND256 : process(INTERP775, INTERP752)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP775 and INTERP752);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP774 <= val after tpd_hl;
            when '1' =>
                INTERP774 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND257 : process(INTERP777, INTERP756)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP777 and INTERP756);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP776 <= val after tpd_hl;
            when '1' =>
                INTERP776 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND258 : process(INTERP779, INTERP760)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP779 and INTERP760);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP778 <= val after tpd_hl;
            when '1' =>
                INTERP778 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND259 : process(INTERP781, INTERP764)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP781 and INTERP764);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP780 <= val after tpd_hl;
            when '1' =>
                INTERP780 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND260 : process(INTERP783, INTERP768)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP783 and INTERP768);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP782 <= val after tpd_hl;
            when '1' =>
                INTERP782 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND261 : process(INTERP785, INTERP772)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP785 and INTERP772);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP784 <= val after tpd_hl;
            when '1' =>
                INTERP784 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND262 : process(INTERP750, INTERP774)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP750 and INTERP774);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP786 <= val after tpd_hl;
            when '1' =>
                INTERP786 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND263 : process(INTERP754, INTERP776)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP754 and INTERP776);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP787 <= val after tpd_hl;
            when '1' =>
                INTERP787 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND264 : process(INTERP758, INTERP778)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP758 and INTERP778);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP788 <= val after tpd_hl;
            when '1' =>
                INTERP788 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND265 : process(INTERP762, INTERP780)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP762 and INTERP780);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP789 <= val after tpd_hl;
            when '1' =>
                INTERP789 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND266 : process(INTERP766, INTERP782)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP766 and INTERP782);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP790 <= val after tpd_hl;
            when '1' =>
                INTERP790 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND267 : process(INTERP770, INTERP784)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP770 and INTERP784);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP791 <= val after tpd_hl;
            when '1' =>
                INTERP791 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV244 : process(INTERP786)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP786);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP792 <= val after tpd_hl;
            when '1' =>
                INTERP792 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV245 : process(INTERP788)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP788);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP793 <= val after tpd_hl;
            when '1' =>
                INTERP793 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV246 : process(INTERP790)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP790);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP794 <= val after tpd_hl;
            when '1' =>
                INTERP794 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV247 : process(INTERP787)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP787);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP795 <= val after tpd_hl;
            when '1' =>
                INTERP795 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV248 : process(INTERP789)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP789);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP796 <= val after tpd_hl;
            when '1' =>
                INTERP796 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND17 : process(INTERP798, INTERP789)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP798 and INTERP789;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP797 <= val after tpd_hl;
            when '1' =>
                INTERP797 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV249 : process(INTERP791)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP791);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP799 <= val after tpd_hl;
            when '1' =>
                INTERP799 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND18 : process(INTERP801, INTERP791)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP801 and INTERP791;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP800 <= val after tpd_hl;
            when '1' =>
                INTERP800 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


 INTERP802 <= not(INTERP735 and INTERP702 and INTERP729 and INTERP792 and INTERP119 and INTERP794 and INTERP793 
             and INTERP120) after tpd_hl;


      AND19 : process(INTERP741, INTERP795)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP741 and INTERP795;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP803 <= val after tpd_hl;
            when '1' =>
                INTERP803 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND20 : process(INTERP805, INTERP795)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP805 and INTERP795;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP804 <= val after tpd_hl;
            when '1' =>
                INTERP804 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND21 : process(INTERP741, INTERP807)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP741 and INTERP807;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP806 <= val after tpd_hl;
            when '1' =>
                INTERP806 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND22 : process(INTERP809, INTERP810)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP809 and INTERP810;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP808 <= val after tpd_hl;
            when '1' =>
                INTERP808 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


 INTERP811 <= INTERP33 and INTERP802 and INTERP31 and INTERP31 after tpd_hl;


      AND24 : process(INTERP259, INTERP796)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP259 and INTERP796;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP812 <= val after tpd_hl;
            when '1' =>
                INTERP812 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND25 : process(INTERP814, INTERP796)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP814 and INTERP796;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP813 <= val after tpd_hl;
            when '1' =>
                INTERP813 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND26 : process(INTERP260, INTERP799)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP260 and INTERP799;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP815 <= val after tpd_hl;
            when '1' =>
                INTERP815 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND27 : process(INTERP817, INTERP799)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP817 and INTERP799;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP816 <= val after tpd_hl;
            when '1' =>
                INTERP816 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


 INTERP818 <= not(INTERP819 and INTERP820 and INTERP806 and INTERP742 and INTERP261) after tpd_hl;


 INTERP821 <= not(INTERP822 and INTERP823 and INTERP803 and INTERP745 and INTERP261) after tpd_hl;


 INTERP824 <= not(INTERP825 and INTERP826 and INTERP803 and INTERP743 and INTERP261) after tpd_hl;


 INTERP827 <= not(INTERP828 and INTERP829 and INTERP804 and INTERP742 and INTERP261) after tpd_hl;


 INTERP830 <= not(INTERP831 and INTERP832 and INTERP808 and INTERP743 and INTERP262) after tpd_hl;


 INTERP833 <= not(INTERP834 and INTERP835 and INTERP806 and INTERP747 and INTERP262) after tpd_hl;


 INTERP836 <= not(INTERP837 and INTERP838 and INTERP808 and INTERP745 and INTERP262) after tpd_hl;


 INTERP839 <= INTERP840 and INTERP841 and INTERP806 and INTERP742 and INTERP261 after tpd_hl;


 INTERP842 <= INTERP843 and INTERP844 and INTERP803 and INTERP745 and INTERP261 after tpd_hl;


 INTERP845 <= INTERP846 and INTERP847 and INTERP803 and INTERP743 and INTERP261 after tpd_hl;


 INTERP848 <= INTERP849 and INTERP850 and INTERP804 and INTERP742 and INTERP261 after tpd_hl;


 INTERP851 <= INTERP852 and INTERP853 and INTERP808 and INTERP743 and INTERP262 after tpd_hl;


 INTERP854 <= INTERP855 and INTERP856 and INTERP806 and INTERP747 and INTERP262 after tpd_hl;


 INTERP857 <= INTERP858 and INTERP859 and INTERP808 and INTERP745 and INTERP262 after tpd_hl;


 INTERP860 <= not(INTERP861 and INTERP816 and INTERP806 and INTERP745 and INTERP261) after tpd_hl;


 INTERP862 <= not(INTERP863 and INTERP816 and INTERP806 and INTERP743 and INTERP261) after tpd_hl;


 INTERP864 <= not(INTERP865 and INTERP816 and INTERP808 and INTERP742 and INTERP261) after tpd_hl;


 INTERP866 <= not(INTERP867 and INTERP816 and INTERP803 and INTERP747 and INTERP261) after tpd_hl;


 INTERP868 <= not(INTERP869 and INTERP816 and INTERP804 and INTERP745 and INTERP262) after tpd_hl;


 INTERP870 <= not(INTERP813 and INTERP871 and INTERP806 and INTERP745 and INTERP262) after tpd_hl;


 INTERP872 <= not(INTERP813 and INTERP873 and INTERP806 and INTERP743 and INTERP262) after tpd_hl;


 INTERP874 <= not(INTERP813 and INTERP875 and INTERP808 and INTERP742 and INTERP262) after tpd_hl;


 INTERP876 <= not(INTERP813 and INTERP877 and INTERP804 and INTERP745 and INTERP262) after tpd_hl;


 INTERP878 <= not(INTERP879 and INTERP816 and INTERP803 and INTERP742 and INTERP147) after tpd_hl;


 INTERP880 <= not(INTERP813 and INTERP881 and INTERP803 and INTERP742 and INTERP147) after tpd_hl;


 INTERP882 <= not(INTERP813 and INTERP816 and INTERP806 and INTERP742 and INTERP147) after tpd_hl;


 INTERP883 <= not(INTERP813 and INTERP816 and INTERP803 and INTERP745 and INTERP147) after tpd_hl;


 INTERP884 <= not(INTERP813 and INTERP816 and INTERP803 and INTERP743 and INTERP147) after tpd_hl;


 INTERP885 <= not(INTERP813 and INTERP816 and INTERP804 and INTERP742 and INTERP147) after tpd_hl;


 INTERP886 <= not(INTERP813 and INTERP815 and INTERP803 and INTERP742 and INTERP147) after tpd_hl;


 INTERP887 <= not(INTERP812 and INTERP816 and INTERP803 and INTERP742 and INTERP147) after tpd_hl;


 INTERP888 <= INTERP889 and INTERP816 and INTERP806 and INTERP745 and INTERP261 after tpd_hl;


 INTERP890 <= INTERP891 and INTERP816 and INTERP806 and INTERP743 and INTERP261 after tpd_hl;


 INTERP892 <= INTERP893 and INTERP816 and INTERP808 and INTERP742 and INTERP261 after tpd_hl;


 INTERP894 <= INTERP895 and INTERP816 and INTERP803 and INTERP747 and INTERP261 after tpd_hl;


 INTERP896 <= INTERP897 and INTERP816 and INTERP804 and INTERP745 and INTERP262 after tpd_hl;


 INTERP898 <= INTERP813 and INTERP899 and INTERP806 and INTERP745 and INTERP262 after tpd_hl;


 INTERP900 <= INTERP813 and INTERP901 and INTERP806 and INTERP743 and INTERP262 after tpd_hl;


 INTERP902 <= INTERP813 and INTERP903 and INTERP808 and INTERP742 and INTERP262 after tpd_hl;


 INTERP904 <= INTERP813 and INTERP905 and INTERP804 and INTERP745 and INTERP262 after tpd_hl;


      NAND293 : process(INTERP839, INTERP34)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP839 and INTERP34);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP906 <= val after tpd_hl;
            when '1' =>
                INTERP906 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV250 : process(INTERP839)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP839);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP907 <= val after tpd_hl;
            when '1' =>
                INTERP907 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND294 : process(INTERP842, INTERP36)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP842 and INTERP36);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP908 <= val after tpd_hl;
            when '1' =>
                INTERP908 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV251 : process(INTERP842)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP842);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP909 <= val after tpd_hl;
            when '1' =>
                INTERP909 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND295 : process(INTERP845, INTERP38)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP845 and INTERP38);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP910 <= val after tpd_hl;
            when '1' =>
                INTERP910 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV252 : process(INTERP845)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP845);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP911 <= val after tpd_hl;
            when '1' =>
                INTERP911 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND296 : process(INTERP848, INTERP40)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP848 and INTERP40);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP912 <= val after tpd_hl;
            when '1' =>
                INTERP912 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV253 : process(INTERP848)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP848);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP913 <= val after tpd_hl;
            when '1' =>
                INTERP913 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND297 : process(INTERP851, INTERP52)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP851 and INTERP52);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP914 <= val after tpd_hl;
            when '1' =>
                INTERP914 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV254 : process(INTERP851)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP851);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP915 <= val after tpd_hl;
            when '1' =>
                INTERP915 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND298 : process(INTERP854, INTERP62)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP854 and INTERP62);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP916 <= val after tpd_hl;
            when '1' =>
                INTERP916 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV255 : process(INTERP854)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP854);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP917 <= val after tpd_hl;
            when '1' =>
                INTERP917 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND299 : process(INTERP857, INTERP64)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP857 and INTERP64);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP918 <= val after tpd_hl;
            when '1' =>
                INTERP918 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV256 : process(INTERP857)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP857);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP919 <= val after tpd_hl;
            when '1' =>
                INTERP919 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


 INTERP920 <= INTERP878 and INTERP880 and INTERP882 and INTERP883 and INTERP884 and INTERP885 and INTERP886
         and INTERP887 after tpd_hl;


      NAND300 : process(INTERP922, INTERP907)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP922 and INTERP907);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP921 <= val after tpd_hl;
            when '1' =>
                INTERP921 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND301 : process(INTERP924, INTERP909)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP924 and INTERP909);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP923 <= val after tpd_hl;
            when '1' =>
                INTERP923 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND302 : process(INTERP926, INTERP911)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP926 and INTERP911);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP925 <= val after tpd_hl;
            when '1' =>
                INTERP925 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND303 : process(INTERP928, INTERP913)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP928 and INTERP913);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP927 <= val after tpd_hl;
            when '1' =>
                INTERP927 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND304 : process(INTERP888, INTERP42)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP888 and INTERP42);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP929 <= val after tpd_hl;
            when '1' =>
                INTERP929 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV257 : process(INTERP888)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP888);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP930 <= val after tpd_hl;
            when '1' =>
                INTERP930 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND305 : process(INTERP890, INTERP44)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP890 and INTERP44);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP931 <= val after tpd_hl;
            when '1' =>
                INTERP931 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV258 : process(INTERP890)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP890);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP932 <= val after tpd_hl;
            when '1' =>
                INTERP932 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND306 : process(INTERP892, INTERP46)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP892 and INTERP46);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP933 <= val after tpd_hl;
            when '1' =>
                INTERP933 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV259 : process(INTERP892)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP892);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP934 <= val after tpd_hl;
            when '1' =>
                INTERP934 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND307 : process(INTERP894, INTERP48)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP894 and INTERP48);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP935 <= val after tpd_hl;
            when '1' =>
                INTERP935 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV260 : process(INTERP894)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP894);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP936 <= val after tpd_hl;
            when '1' =>
                INTERP936 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND308 : process(INTERP896, INTERP50)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP896 and INTERP50);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP937 <= val after tpd_hl;
            when '1' =>
                INTERP937 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV261 : process(INTERP896)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP896);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP938 <= val after tpd_hl;
            when '1' =>
                INTERP938 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND309 : process(INTERP940, INTERP915)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP940 and INTERP915);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP939 <= val after tpd_hl;
            when '1' =>
                INTERP939 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND310 : process(INTERP898, INTERP54)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP898 and INTERP54);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP941 <= val after tpd_hl;
            when '1' =>
                INTERP941 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV262 : process(INTERP898)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP898);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP942 <= val after tpd_hl;
            when '1' =>
                INTERP942 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND311 : process(INTERP900, INTERP56)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP900 and INTERP56);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP943 <= val after tpd_hl;
            when '1' =>
                INTERP943 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV263 : process(INTERP900)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP900);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP944 <= val after tpd_hl;
            when '1' =>
                INTERP944 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND312 : process(INTERP902, INTERP58)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP902 and INTERP58);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP945 <= val after tpd_hl;
            when '1' =>
                INTERP945 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV264 : process(INTERP902)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP902);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP946 <= val after tpd_hl;
            when '1' =>
                INTERP946 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND313 : process(INTERP904, INTERP60)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP904 and INTERP60);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP947 <= val after tpd_hl;
            when '1' =>
                INTERP947 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV265 : process(INTERP904)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP904);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP948 <= val after tpd_hl;
            when '1' =>
                INTERP948 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND314 : process(INTERP950, INTERP917)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP950 and INTERP917);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP949 <= val after tpd_hl;
            when '1' =>
                INTERP949 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND315 : process(INTERP952, INTERP919)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP952 and INTERP919);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP951 <= val after tpd_hl;
            when '1' =>
                INTERP951 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


 INTERP953 <= not(INTERP818 and INTERP821 and INTERP824 and INTERP827 and INTERP860 and INTERP862 and INTERP864 
             and INTERP866) after tpd_hl;


 INTERP954 <= not(INTERP868 and INTERP830 and INTERP870 and INTERP872 and INTERP874 and INTERP876 and INTERP833 
             and INTERP836) after tpd_hl;


 INTERP955 <= INTERP818 and INTERP821 and INTERP824 and INTERP827 and INTERP860 and INTERP862 and INTERP864
         and INTERP866 after tpd_hl;


 INTERP956 <= INTERP868 and INTERP830 and INTERP870 and INTERP872 and INTERP874 and INTERP876 and INTERP833
         and INTERP836 after tpd_hl;


      NAND318 : process(INTERP906, INTERP921)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP906 and INTERP921);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(0) <= val after tpd_hl;
            when '1' =>
                OUTPI(0) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND319 : process(INTERP908, INTERP923)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP908 and INTERP923);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(1) <= val after tpd_hl;
            when '1' =>
                OUTPI(1) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND320 : process(INTERP910, INTERP925)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP910 and INTERP925);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(2) <= val after tpd_hl;
            when '1' =>
                OUTPI(2) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND321 : process(INTERP912, INTERP927)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP912 and INTERP927);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(3) <= val after tpd_hl;
            when '1' =>
                OUTPI(3) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND322 : process(INTERP958, INTERP930)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP958 and INTERP930);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP957 <= val after tpd_hl;
            when '1' =>
                INTERP957 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND323 : process(INTERP960, INTERP932)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP960 and INTERP932);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP959 <= val after tpd_hl;
            when '1' =>
                INTERP959 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND324 : process(INTERP962, INTERP934)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP962 and INTERP934);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP961 <= val after tpd_hl;
            when '1' =>
                INTERP961 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND325 : process(INTERP964, INTERP936)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP964 and INTERP936);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP963 <= val after tpd_hl;
            when '1' =>
                INTERP963 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND326 : process(INTERP966, INTERP938)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP966 and INTERP938);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP965 <= val after tpd_hl;
            when '1' =>
                INTERP965 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND327 : process(INTERP914, INTERP939)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP914 and INTERP939);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(4) <= val after tpd_hl;
            when '1' =>
                OUTPI(4) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND328 : process(INTERP968, INTERP942)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP968 and INTERP942);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP967 <= val after tpd_hl;
            when '1' =>
                INTERP967 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND329 : process(INTERP970, INTERP944)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP970 and INTERP944);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP969 <= val after tpd_hl;
            when '1' =>
                INTERP969 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND330 : process(INTERP972, INTERP946)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP972 and INTERP946);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP971 <= val after tpd_hl;
            when '1' =>
                INTERP971 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND331 : process(INTERP974, INTERP948)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP974 and INTERP948);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP973 <= val after tpd_hl;
            when '1' =>
                INTERP973 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND332 : process(INTERP916, INTERP949)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP916 and INTERP949);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(5) <= val after tpd_hl;
            when '1' =>
                OUTPI(5) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND333 : process(INTERP918, INTERP951)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP918 and INTERP951);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(6) <= val after tpd_hl;
            when '1' =>
                OUTPI(6) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND47 : process(INTERP953, INTERP24)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP953 and INTERP24;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP975 <= val after tpd_hl;
            when '1' =>
                INTERP975 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND48 : process(INTERP954, INTERP25)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP954 and INTERP25;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP976 <= val after tpd_hl;
            when '1' =>
                INTERP976 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND334 : process(INTERP929, INTERP957)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP929 and INTERP957);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(7) <= val after tpd_hl;
            when '1' =>
                OUTPI(7) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND335 : process(INTERP931, INTERP959)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP931 and INTERP959);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(8) <= val after tpd_hl;
            when '1' =>
                OUTPI(8) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND336 : process(INTERP933, INTERP961)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP933 and INTERP961);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(9) <= val after tpd_hl;
            when '1' =>
                OUTPI(9) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND337 : process(INTERP935, INTERP963)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP935 and INTERP963);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(10) <= val after tpd_hl;
            when '1' =>
                OUTPI(10) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND338 : process(INTERP937, INTERP965)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP937 and INTERP965);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(11) <= val after tpd_hl;
            when '1' =>
                OUTPI(11) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND339 : process(INTERP941, INTERP967)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP941 and INTERP967);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(12) <= val after tpd_hl;
            when '1' =>
                OUTPI(12) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND340 : process(INTERP943, INTERP969)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP943 and INTERP969);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(13) <= val after tpd_hl;
            when '1' =>
                OUTPI(13) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND341 : process(INTERP945, INTERP971)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP945 and INTERP971);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(14) <= val after tpd_hl;
            when '1' =>
                OUTPI(14) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND342 : process(INTERP947, INTERP973)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP947 and INTERP973);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(15) <= val after tpd_hl;
            when '1' =>
                OUTPI(15) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND343 : process(INTERP955, INTERP956)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP955 and INTERP956);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP978 <= val after tpd_hl;
            when '1' =>
                INTERP978 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


 INTERP979 <= INTERP33 and INTERP802 and INP(31) and INTERP977 after tpd_hl;


      NAND344 : process(INTERP975, INTERP709)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP975 and INTERP709);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP980 <= val after tpd_hl;
            when '1' =>
                INTERP980 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV266 : process(INTERP975)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP975);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP981 <= val after tpd_hl;
            when '1' =>
                INTERP981 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND345 : process(INTERP976, INTERP710)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP976 and INTERP710);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP982 <= val after tpd_hl;
            when '1' =>
                INTERP982 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV267 : process(INTERP976)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP976);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP983 <= val after tpd_hl;
            when '1' =>
                INTERP983 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NOR0 : process(INTERP811, INTERP979)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP811 or INTERP979);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(16) <= val after tpd_hl;
            when '1' =>
                OUTPI(16) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND346 : process(INTERP670, INTERP981)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP670 and INTERP981);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP994 <= val after tpd_hl;
            when '1' =>
                INTERP994 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND347 : process(INTERP671, INTERP983)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP671 and INTERP983);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP995 <= val after tpd_hl;
            when '1' =>
                INTERP995 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND348 : process(INTERP980, INTERP994)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP980 and INTERP994);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP998 <= val after tpd_hl;
            when '1' =>
                INTERP998 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND349 : process(INTERP982, INTERP995)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP982 and INTERP995);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP999 <= val after tpd_hl;
            when '1' =>
                INTERP999 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND350 : process(INTERP984, INTERP737)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP984 and INTERP737);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1000 <= val after tpd_hl;
            when '1' =>
                INTERP1000 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND351 : process(INTERP986, INTERP738)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP986 and INTERP738);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1001 <= val after tpd_hl;
            when '1' =>
                INTERP1001 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND352 : process(INTERP988, INTERP646)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP988 and INTERP646);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1002 <= val after tpd_hl;
            when '1' =>
                INTERP1002 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND353 : process(INTERP990, INTERP622)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP990 and INTERP622);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1003 <= val after tpd_hl;
            when '1' =>
                INTERP1003 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND354 : process(INTERP992, INTERP662)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP992 and INTERP662);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1004 <= val after tpd_hl;
            when '1' =>
                INTERP1004 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV268 : process(INTERP984)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP984);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1005 <= val after tpd_hl;
            when '1' =>
                INTERP1005 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV269 : process(INTERP986)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP986);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1006 <= val after tpd_hl;
            when '1' =>
                INTERP1006 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV270 : process(INTERP988)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP988);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1007 <= val after tpd_hl;
            when '1' =>
                INTERP1007 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV271 : process(INTERP990)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP990);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1008 <= val after tpd_hl;
            when '1' =>
                INTERP1008 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV272 : process(INTERP992)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP992);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1009 <= val after tpd_hl;
            when '1' =>
                INTERP1009 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV273 : process(INTERP996)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP996);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1010 <= val after tpd_hl;
            when '1' =>
                INTERP1010 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND355 : process(INTERP996, INTERP682)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP996 and INTERP682);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1011 <= val after tpd_hl;
            when '1' =>
                INTERP1011 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND356 : process(INTERP730, INTERP1005)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP730 and INTERP1005);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1012 <= val after tpd_hl;
            when '1' =>
                INTERP1012 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND357 : process(INTERP731, INTERP1006)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP731 and INTERP1006);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1013 <= val after tpd_hl;
            when '1' =>
                INTERP1013 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND358 : process(INTERP1015, INTERP1007)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP1015 and INTERP1007);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1014 <= val after tpd_hl;
            when '1' =>
                INTERP1014 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND359 : process(INTERP1017, INTERP1008)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP1017 and INTERP1008);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1016 <= val after tpd_hl;
            when '1' =>
                INTERP1016 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND360 : process(INTERP1019, INTERP1009)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP1019 and INTERP1009);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1018 <= val after tpd_hl;
            when '1' =>
                INTERP1018 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND361 : process(INTERP998, INTERP99)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP998 and INTERP99);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1020 <= val after tpd_hl;
            when '1' =>
                INTERP1020 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV274 : process(INTERP998)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP998);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1021 <= val after tpd_hl;
            when '1' =>
                INTERP1021 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND362 : process(INTERP999, INTERP100)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP999 and INTERP100);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1022 <= val after tpd_hl;
            when '1' =>
                INTERP1022 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV275 : process(INTERP999)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP999);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1023 <= val after tpd_hl;
            when '1' =>
                INTERP1023 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND363 : process(INTERP659, INTERP1010)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP659 and INTERP1010);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1024 <= val after tpd_hl;
            when '1' =>
                INTERP1024 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND364 : process(INTERP1012, INTERP1000)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP1012 and INTERP1000);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1025 <= val after tpd_hl;
            when '1' =>
                INTERP1025 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND365 : process(INTERP1013, INTERP1001)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP1013 and INTERP1001);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1026 <= val after tpd_hl;
            when '1' =>
                INTERP1026 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND366 : process(INTERP1014, INTERP1002)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP1014 and INTERP1002);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1027 <= val after tpd_hl;
            when '1' =>
                INTERP1027 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND367 : process(INTERP1016, INTERP1003)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP1016 and INTERP1003);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1028 <= val after tpd_hl;
            when '1' =>
                INTERP1028 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND368 : process(INTERP1018, INTERP1004)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP1018 and INTERP1004);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1029 <= val after tpd_hl;
            when '1' =>
                INTERP1029 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND369 : process(INTERP94, INTERP1021)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP94 and INTERP1021);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1030 <= val after tpd_hl;
            when '1' =>
                INTERP1030 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND370 : process(INTERP96, INTERP1023)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP96 and INTERP1023);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1031 <= val after tpd_hl;
            when '1' =>
                INTERP1031 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND371 : process(INTERP1024, INTERP1011)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP1024 and INTERP1011);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1032 <= val after tpd_hl;
            when '1' =>
                INTERP1032 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND57 : process(INTERP1025, INTERP66)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP1025 and INTERP66;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(17) <= val after tpd_hl;
            when '1' =>
                OUTPI(17) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND58 : process(INTERP68, INTERP1026)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP68 and INTERP1026;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(18) <= val after tpd_hl;
            when '1' =>
                OUTPI(18) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND59 : process(INTERP72, INTERP1027)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP72 and INTERP1027;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(19) <= val after tpd_hl;
            when '1' =>
                OUTPI(19) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND60 : process(INTERP1028, INTERP74)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP1028 and INTERP74;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(20) <= val after tpd_hl;
            when '1' =>
                OUTPI(20) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND61 : process(INTERP76, INTERP1029)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP76 and INTERP1029;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(21) <= val after tpd_hl;
            when '1' =>
                OUTPI(21) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND372 : process(INTERP1020, INTERP1030)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP1020 and INTERP1030);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(22) <= val after tpd_hl;
            when '1' =>
                OUTPI(22) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND373 : process(INTERP1022, INTERP1031)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP1022 and INTERP1031);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(23) <= val after tpd_hl;
            when '1' =>
                OUTPI(23) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND374 : process(INTERP1032, INTERP424)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP1032 and INTERP424);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1033 <= val after tpd_hl;
            when '1' =>
                INTERP1033 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      INV276 : process(INTERP1032)
        variable val,ex_value : bit := '0';

    begin
        val := not(INTERP1032);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1034 <= val after tpd_hl;
            when '1' =>
                INTERP1034 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND375 : process(INTERP384, INTERP1034)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP384 and INTERP1034);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1035 <= val after tpd_hl;
            when '1' =>
                INTERP1035 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      NAND376 : process(INTERP1033, INTERP1035)
        variable val,ex_value : bit := '0';
    begin
        val := not(INTERP1033 and INTERP1035);

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                INTERP1036 <= val after tpd_hl;
            when '1' =>
                INTERP1036 <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;


      AND62 : process(INTERP1036, INTERP70)
        variable val,ex_value : bit := '0';
    begin
        val := INTERP1036 and INTERP70;

        if val /= ex_value then
          ex_value := val;
          case val is 
            when '0' =>
                OUTPI(24) <= val after tpd_hl;
            when '1' =>
                OUTPI(24) <= val after tpd_lh;
            when others =>
          end case;
        end if;  
    end process;

  BUFFER_OUT : OUTP <= OUTPI;

p:process

 file test_in : text is in "iscas5.in";
 variable L : line;
 variable x : bit_vector(0 to 32);
 variable y : bit;
 begin
  while(not(endfile(test_in))) loop
   readline(test_in,L);
   read(L,x);
   read(L,y);
   INP <= x;
   H <= y; 
   wait for 200 fs;
 end loop;
 wait;
end process;

printout:process
 variable outline : LINE;
 variable S1 : string(1 to 6) := " I1 = ";
 variable S2 : string(1 to 6) := " I2 = ";
 variable S3 : string(1 to 5) := "OP = ";
 file outfile: TEXT is out "ISCAS85_5.out";

begin
 wait for 200 fs;
 write(outline, now);
 writeline(outfile,outline);
 write(outline,S1);
 write(outline,INP);
 write(outline,S2);
 write(outline,H);
 writeline(outfile,outline);
 write(outline,S3);
 write(outline,OUTP);
 writeline(outfile,outline);
 wait on INP,H ;
end process;

end DEMO;



